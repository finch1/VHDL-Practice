--enc_int