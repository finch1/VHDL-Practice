//Legal Notice: (C)2008 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module dut (
             // inputs:
              asi_sink_data,
              csi_clock_clk,
              csi_clock_reset,

             // outputs:
              aso_source_data
           )
;

  output  [ 15: 0] aso_source_data;
  input   [ 15: 0] asi_sink_data;
  input            csi_clock_clk;
  input            csi_clock_reset;

  wire    [ 15: 0] aso_source_data;
  my_dut the_my_dut
    (
      .asi_sink_data   (asi_sink_data),
      .aso_source_data (aso_source_data),
      .csi_clock_clk   (csi_clock_clk),
      .csi_clock_reset (csi_clock_reset)
    );


endmodule

