-- megafunction wizard: %altasmi_parallel%
-- generation: standard
-- version: wm1.0
-- module: altasmi_parallel 

-- ============================================================
-- file name: altasmi.vhd
-- megafunction name(s):
-- 			altasmi_parallel
--
-- simulation library files(s):
-- 			
-- ============================================================
-- ************************************************************
-- this is a wizard-generated file. do not edit this file!
--
-- 13.1.0 build 162 10/23/2013 sj web edition
-- ************************************************************


--copyright (c) 1991-2013 altera corporation
--your use of altera corporation's design tools, logic functions 
--and other software and tools, and its ampp partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the altera program license 
--subscription agreement, altera megacore function license 
--agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by altera and sold by 
--altera or its authorized distributors.  please refer to the 
--applicable agreement for further details.


--altasmi_parallel cbx_auto_blackbox="all" data_width="standard" device_family="cyclone iii" epcs_type="epcs4" page_size=1 port_bulk_erase="port_unused" port_die_erase="port_unused" port_en4b_addr="port_unused" port_ex4b_addr="port_unused" port_fast_read="port_unused" port_illegal_erase="port_unused" port_illegal_write="port_used" port_rdid_out="port_unused" port_read_address="port_unused" port_read_dummyclk="port_unused" port_read_rdid="port_unused" port_read_sid="port_unused" port_read_status="port_unused" port_sector_erase="port_unused" port_sector_protect="port_unused" port_shift_bytes="port_unused" port_wren="port_used" port_write="port_used" use_asmiblock="on" use_eab="on" write_dummy_clk=0 addr busy clkin data_valid datain dataout illegal_write rden read reset wren write intended_device_family="cyclone iii" altera_internal_options=suppress_da_rule_internal=c106
--version_begin 13.1 cbx_a_gray2bin 2013:10:24:09:15:20:sj cbx_a_graycounter 2013:10:24:09:15:20:sj cbx_altasmi_parallel 2013:10:24:09:15:20:sj cbx_altdpram 2013:10:24:09:15:20:sj cbx_altsyncram 2013:10:24:09:15:20:sj cbx_arriav 2013:10:24:09:15:20:sj cbx_cyclone 2013:10:24:09:15:20:sj cbx_cycloneii 2013:10:24:09:15:20:sj cbx_fifo_common 2013:10:24:09:15:20:sj cbx_lpm_add_sub 2013:10:24:09:15:20:sj cbx_lpm_compare 2013:10:24:09:15:20:sj cbx_lpm_counter 2013:10:24:09:15:20:sj cbx_lpm_decode 2013:10:24:09:15:20:sj cbx_lpm_mux 2013:10:24:09:15:20:sj cbx_mgl 2013:10:24:09:16:30:sj cbx_nightfury 2013:10:24:09:15:19:sj cbx_scfifo 2013:10:24:09:15:20:sj cbx_stratix 2013:10:24:09:15:20:sj cbx_stratixii 2013:10:24:09:15:20:sj cbx_stratixiii 2013:10:24:09:15:20:sj cbx_stratixv 2013:10:24:09:15:20:sj cbx_util_mgl 2013:10:24:09:15:20:sj  version_end

 library altera_mf;
 use altera_mf.all;

 library cycloneii;
 use cycloneii.all;

--synthesis_resources = a_graycounter 4 cycloneii_asmiblock 1 lut 27 mux21 1 reg 96 
 library ieee;
 use ieee.std_logic_1164.all;

 entity  altasmi_altasmi_parallel_3kj2 is 
	 port 
	 ( 
		 addr	:	in  std_logic_vector (23 downto 0);
		 busy	:	out  std_logic;
		 clkin	:	in  std_logic;
		 data_valid	:	out  std_logic;
		 datain	:	in  std_logic_vector (7 downto 0) := (others => '0');
		 dataout	:	out  std_logic_vector (7 downto 0);
		 illegal_write	:	out  std_logic;
		 rden	:	in  std_logic;
		 read	:	in  std_logic := '0';
		 reset	:	in  std_logic := '0';
		 wren	:	in  std_logic := '1';
		 write	:	in  std_logic := '0'
	 ); 
 end altasmi_altasmi_parallel_3kj2;

 architecture rtl of altasmi_altasmi_parallel_3kj2 is

	 attribute synthesis_clearbox : natural;
	 attribute synthesis_clearbox of rtl : architecture is 2;
	 attribute altera_attribute : string;
	 attribute altera_attribute of rtl : architecture is "suppress_da_rule_internal=c106";

	 signal  wire_addbyte_cntr_w_lg_w_q_range158w163w	:	std_logic_vector (0 downto 0);
	 signal  wire_addbyte_cntr_w_lg_w_q_range161w162w	:	std_logic_vector (0 downto 0);
	 signal  wire_addbyte_cntr_clk_en	:	std_logic;
	 signal  wire_stage_cntr_w157w	:	std_logic_vector (0 downto 0);
	 signal  wire_addbyte_cntr_clock	:	std_logic;
	 signal  wire_addbyte_cntr_q	:	std_logic_vector (2 downto 0);
	 signal  wire_addbyte_cntr_sclr	:	std_logic;
	 signal  wire_w_lg_end_operation100w	:	std_logic_vector (0 downto 0);
	 signal  wire_addbyte_cntr_w_q_range161w	:	std_logic_vector (0 downto 0);
	 signal  wire_addbyte_cntr_w_q_range158w	:	std_logic_vector (0 downto 0);
	 signal  wire_gen_cntr_w_lg_w_q_range113w114w	:	std_logic_vector (0 downto 0);
	 signal  wire_gen_cntr_w_lg_w_q_range111w112w	:	std_logic_vector (0 downto 0);
	 signal  wire_gen_cntr_clk_en	:	std_logic;
	 signal  wire_w_lg_w_lg_w_lg_in_operation40w41w42w	:	std_logic_vector (0 downto 0);
	 signal  wire_gen_cntr_q	:	std_logic_vector (2 downto 0);
	 signal  wire_gen_cntr_sclr	:	std_logic;
	 signal  wire_w_lg_w_lg_end1_cyc_reg_in_wire43w44w	:	std_logic_vector (0 downto 0);
	 signal  wire_gen_cntr_w_q_range111w	:	std_logic_vector (0 downto 0);
	 signal  wire_gen_cntr_w_q_range113w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w332w333w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w332w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w337w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range103w106w329w330w331w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range103w106w334w335w336w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range103w104w105w343w344w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range103w108w420w421w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range103w106w329w330w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range103w106w354w355w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range103w106w334w335w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range103w104w105w343w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_lg_w_q_range103w108w420w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_lg_w_q_range103w106w329w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_lg_w_q_range103w106w354w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_lg_w_q_range103w106w334w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_lg_w_q_range103w106w154w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_lg_w_q_range103w106w327w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range102w107w133w134w135w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_lg_w_q_range102w107w133w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_lg_w_q_range103w104w105w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_q_range103w108w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_q_range103w106w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range102w107w133w134w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_q_range102w107w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_lg_w_q_range103w104w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_clk_en	:	std_logic;
	 signal  wire_w_lg_w_lg_w_lg_w96w97w98w99w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_q	:	std_logic_vector (1 downto 0);
	 signal  wire_stage_cntr_sclr	:	std_logic;
	 signal  wire_stage_cntr_w_q_range102w	:	std_logic_vector (0 downto 0);
	 signal  wire_stage_cntr_w_q_range103w	:	std_logic_vector (0 downto 0);
	 signal  wire_wrstage_cntr_w_lg_w_q_range524w525w	:	std_logic_vector (0 downto 0);
	 signal  wire_wrstage_cntr_w_lg_w_q_range522w523w	:	std_logic_vector (0 downto 0);
	 signal  wire_wrstage_cntr_clk_en	:	std_logic;
	 signal  wire_w_lg_w_lg_w_lg_w_lg_w517w518w519w520w521w	:	std_logic_vector (0 downto 0);
	 signal  wire_wrstage_cntr_clock	:	std_logic;
	 signal  wire_wrstage_cntr_q	:	std_logic_vector (1 downto 0);
	 signal  wire_wrstage_cntr_w_q_range522w	:	std_logic_vector (0 downto 0);
	 signal  wire_wrstage_cntr_w_q_range524w	:	std_logic_vector (0 downto 0);
	 signal  wire_cycloneii_asmiblock2_data0out	:	std_logic;
	 signal  wire_cycloneii_asmiblock2_sdoin	:	std_logic;
	 signal  wire_w_lg_sdoin_wire320w	:	std_logic_vector (0 downto 0);
	 signal	 add_msb_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 wire_add_msb_reg_ena	:	std_logic;
	 signal	 wire_addr_reg_d	:	std_logic_vector (23 downto 0);
	 signal	 addr_reg	:	std_logic_vector(23 downto 0)
	 -- synopsys translate_off
	  := (others => '0')
	 -- synopsys translate_on
	 ;
	 signal	 wire_addr_reg_ena	:	std_logic_vector(23 downto 0);
	 signal  wire_addr_reg_w_q_range574w	:	std_logic_vector (0 downto 0);
	 signal  wire_addr_reg_w_q_range581w	:	std_logic_vector (0 downto 0);
	 signal  wire_addr_reg_w_q_range393w	:	std_logic_vector (22 downto 0);
	 signal  wire_addr_reg_w_q_range586w	:	std_logic_vector (0 downto 0);
	 signal	 wire_asmi_opcode_reg_d	:	std_logic_vector (7 downto 0);
	 signal	 asmi_opcode_reg	:	std_logic_vector(7 downto 0)
	 -- synopsys translate_off
	  := (others => '0')
	 -- synopsys translate_on
	 ;
	 signal	 wire_asmi_opcode_reg_ena	:	std_logic_vector(7 downto 0);
	 signal  wire_asmi_opcode_reg_w_q_range168w	:	std_logic_vector (6 downto 0);
	 signal	 busy_det_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 clr_read_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 clr_read_reg2	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 clr_rstat_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 clr_write_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 clr_write_reg2	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 wire_datain_reg_d	:	std_logic_vector (7 downto 0);
	 signal	 datain_reg	:	std_logic_vector(7 downto 0)
	 -- synopsys translate_off
	  := (others => '0')
	 -- synopsys translate_on
	 ;
	 signal	 wire_datain_reg_ena	:	std_logic_vector(7 downto 0);
	 signal  wire_datain_reg_w_q_range614w	:	std_logic_vector (6 downto 0);
	 signal	 do_wrmemadd_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 dvalid_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 wire_dvalid_reg_ena	:	std_logic;
	 signal	 wire_dvalid_reg_sclr	:	std_logic;
	 signal	 dvalid_reg2	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 end1_cyc_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 end1_cyc_reg2	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 end_op_hdlyreg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 end_op_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 end_rbyte_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 wire_end_rbyte_reg_ena	:	std_logic;
	 signal	 wire_end_rbyte_reg_sclr	:	std_logic;
	 signal	 end_read_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 ill_write_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 illegal_write_prot_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 ncs_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 wire_ncs_reg_sclr	:	std_logic;
	 signal  wire_ncs_reg_w_lg_q380w	:	std_logic_vector (0 downto 0);
	 signal	 wire_read_data_reg_d	:	std_logic_vector (7 downto 0);
	 signal	 read_data_reg	:	std_logic_vector(7 downto 0)
	 -- synopsys translate_off
	  := (others => '0')
	 -- synopsys translate_on
	 ;
	 signal	 wire_read_data_reg_ena	:	std_logic_vector(7 downto 0);
	 signal	 wire_read_dout_reg_d	:	std_logic_vector (7 downto 0);
	 signal	 read_dout_reg	:	std_logic_vector(7 downto 0)
	 -- synopsys translate_off
	  := (others => '0')
	 -- synopsys translate_on
	 ;
	 signal	 wire_read_dout_reg_ena	:	std_logic_vector(7 downto 0);
	 signal	 read_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 wire_read_reg_ena	:	std_logic;
	 signal	 shift_op_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 stage2_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 stage3_dly_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 stage3_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 stage4_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 start_wrpoll_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 wire_start_wrpoll_reg_ena	:	std_logic;
	 signal	 start_wrpoll_reg2	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 wire_statreg_int_d	:	std_logic_vector (7 downto 0);
	 signal	 statreg_int	:	std_logic_vector(7 downto 0)
	 -- synopsys translate_off
	  := (others => '0')
	 -- synopsys translate_on
	 ;
	 signal	 wire_statreg_int_ena	:	std_logic_vector(7 downto 0);
	 signal	 write_prot_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 wire_write_prot_reg_ena	:	std_logic;
	 signal	 write_prot_reg2	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 write_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 wire_write_reg_ena	:	std_logic;
	 signal	 write_rstat_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	 wrsdoin_reg	:	std_logic
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 signal	wire_mux211_dataout	:	std_logic;
	 signal  wire_w_lg_w_lg_w655w656w657w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w655w656w	:	std_logic_vector (0 downto 0);
	 signal  wire_w287w	:	std_logic_vector (0 downto 0);
	 signal  wire_w227w	:	std_logic_vector (6 downto 0);
	 signal  wire_w285w	:	std_logic_vector (0 downto 0);
	 signal  wire_w220w	:	std_logic_vector (6 downto 0);
	 signal  wire_w655w	:	std_logic_vector (0 downto 0);
	 signal  wire_w477w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_load_opcode184w185w186w271w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_load_opcode184w185w186w187w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_load_opcode189w190w191w273w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_load_opcode189w190w191w192w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_load_opcode223w224w225w226w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_load_opcode194w195w196w275w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_load_opcode194w195w196w197w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_load_opcode235w236w237w293w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_load_opcode235w236w237w238w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_load_opcode216w217w218w219w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_do_read359w360w361w362w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_do_write651w652w653w654w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w530w641w642w658w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_do_read407w474w475w476w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_do_sec_erase54w416w417w418w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_do_write628w629w630w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_load_opcode184w185w186w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_load_opcode189w190w191w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_load_opcode199w204w279w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_load_opcode199w204w205w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_load_opcode199w200w277w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_load_opcode199w200w201w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_load_opcode223w224w225w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_load_opcode194w195w196w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_load_opcode235w236w237w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_load_opcode216w217w218w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_bp2_wire547w548w549w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_bp2_wire547w548w552w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_bp2_wire547w554w555w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_bp2_wire547w554w557w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_do_read359w360w361w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_do_read359w360w419w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_do_write651w652w653w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w530w641w642w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_do_read407w474w475w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_do_sec_erase54w416w417w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_bp2_wire559w560w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_bp2_wire559w562w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_bp2_wire564w565w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_bp2_wire564w567w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_do_4baddr176w177w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_do_ex4baddr171w172w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_do_polling500w501w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_do_read_stat123w124w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_do_write207w208w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_do_write628w629w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_do_write63w338w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode178w267w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode178w179w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode173w265w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode173w174w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode209w281w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode209w210w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode184w185w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode189w190w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode229w289w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode229w230w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode232w291w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode232w233w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode212w283w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode212w213w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode240w295w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode240w241w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode243w297w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode243w244w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode199w204w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode199w200w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode223w224w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode194w195w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode235w236w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode181w269w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode181w182w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_load_opcode216w217w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_stage3_wire45w46w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_start_poll345w346w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_bp2_wire547w548w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_bp2_wire547w554w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_do_read359w360w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_do_write651w652w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w517w518w519w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w530w641w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_do_write72w116w117w516w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_do_write72w116w117w130w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_do_write72w73w408w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_do_read407w474w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_do_read_rdid125w126w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_do_sec_erase54w416w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_end_operation502w503w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_rden_wire412w413w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_addr_overdie402w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_addr_overdie392w	:	std_logic_vector (22 downto 0);
	 signal  wire_w_lg_bp2_wire559w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_bp2_wire564w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_4baddr176w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_bulk_erase339w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_ex4baddr171w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_polling500w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_read_nonvolatile325w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_read_stat123w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_write207w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_write628w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_write70w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_write63w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_load_opcode178w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_load_opcode173w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_load_opcode209w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_load_opcode184w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_load_opcode189w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_load_opcode229w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_load_opcode232w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_load_opcode212w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_load_opcode240w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_load_opcode243w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_load_opcode199w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_load_opcode223w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_load_opcode194w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_load_opcode235w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_load_opcode181w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_load_opcode216w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_not_busy404w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_not_busy396w	:	std_logic_vector (22 downto 0);
	 signal  wire_w_lg_not_busy622w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_not_busy617w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_shift_opcode169w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_stage3_wire410w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_stage3_wire441w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_stage3_wire55w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_stage3_wire45w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_stage3_wire394w	:	std_logic_vector (22 downto 0);
	 signal  wire_w_lg_stage4_wire443w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_stage4_wire411w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_stage4_wire615w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_start_poll345w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_wren_wire631w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_mask_prot_range568w575w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_mask_prot_range571w582w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_mask_prot_range573w587w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_do_write63w357w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w119w120w121w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_addr_overdie490w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_bp0_wire545w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_bp1_wire546w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_bp2_wire547w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_busy_wire1w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_clkin_wire101w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_4baddr647w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_bulk_erase649w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_die_erase648w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_ex4baddr646w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_fast_read358w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_memadd425w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_polling203w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_read359w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_read_rdid51w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_read_stat52w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_read_volatile215w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_sec_erase650w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_wren53w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_write651w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_write_rstat627w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_write_volatile222w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_end_add_cycle83w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_end_fast_read77w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_end_ophdly39w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_end_pgwr_data62w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_end_read80w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_rden_wire492w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_read_rdid_wire9w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_read_sid_wire8w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_sec_protect_wire7w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_st_busy_wire127w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_start_poll122w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_write_prot_true515w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_write_wire17w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_pagewr_buf_not_empty_range68w69w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_w530w641w642w658w659w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_load_opcode243w297w298w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_load_opcode243w244w245w	:	std_logic_vector (6 downto 0);
	 signal  wire_w517w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_do_write72w73w408w409w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_end_operation502w503w504w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_rden_wire412w413w414w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_not_busy404w405w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_not_busy396w397w	:	std_logic_vector (22 downto 0);
	 signal  wire_w_lg_w_lg_not_busy617w618w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_stage4_wire443w444w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_wren_wire631w632w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_load_opcode243w297w298w299w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_load_opcode243w244w245w246w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w517w518w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_rden_wire412w413w414w415w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_not_busy396w397w398w	:	std_logic_vector (22 downto 0);
	 signal  wire_w300w	:	std_logic_vector (0 downto 0);
	 signal  wire_w247w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w300w301w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w247w248w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_w300w301w302w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w247w248w249w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w300w301w302w303w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w247w248w249w250w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_w300w301w302w303w304w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_w247w248w249w250w251w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w300w301w302w303w304w305w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w247w248w249w250w251w252w	:	std_logic_vector (6 downto 0);
	 signal  wire_w306w	:	std_logic_vector (0 downto 0);
	 signal  wire_w253w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w306w307w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w253w254w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_w306w307w308w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w253w254w255w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w306w307w308w309w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w253w254w255w256w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_w306w307w308w309w310w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_w253w254w255w256w257w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w306w307w308w309w310w311w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w253w254w255w256w257w258w	:	std_logic_vector (6 downto 0);
	 signal  wire_w312w	:	std_logic_vector (0 downto 0);
	 signal  wire_w259w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w312w313w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w259w260w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_w259w260w261w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_lg_w_lg_w151w152w153w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w151w152w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w119w120w	:	std_logic_vector (0 downto 0);
	 signal  wire_w151w	:	std_logic_vector (0 downto 0);
	 signal  wire_w530w	:	std_logic_vector (0 downto 0);
	 signal  wire_w119w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_do_read407w428w429w430w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_do_read_sid147w148w149w150w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_do_write72w116w117w529w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_w_lg_do_write72w116w117w118w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_bp3_wire539w540w541w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_do_read407w428w429w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_do_read_sid147w148w149w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_do_read_stat438w439w440w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_do_sec_erase532w533w534w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_lg_do_write72w116w117w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_bp3_wire539w540w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_do_read407w442w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_do_read407w428w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_do_read_sid147w148w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_do_read_stat438w439w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_do_sec_erase532w533w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_do_write72w116w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_do_write72w73w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_lg_w_prot_wire_range551w570w572w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_bp3_wire539w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_data0out_wire446w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_4baddr341w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_ex4baddr340w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_read407w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_read_rdid125w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_read_sid147w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_read_stat438w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_sec_erase54w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_sec_erase532w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_wren342w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_do_write72w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_end_operation502w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_load_opcode315w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_rden_wire412w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_mask_prot_add_range583w597w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_mask_prot_add_range588w601w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_mask_prot_check_range585w595w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_mask_prot_check_range590w599w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_prot_wire_range551w570w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_mask_prot_range568w578w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_mask_prot_range571w584w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_lg_w_mask_prot_range573w589w	:	std_logic_vector (0 downto 0);
	 signal  addr_overdie :	std_logic;
	 signal  addr_overdie_pos :	std_logic;
	 signal  addr_reg_overdie :	std_logic_vector (23 downto 0);
	 signal  b4addr_opcode :	std_logic_vector (7 downto 0);
	 signal  be_write_prot :	std_logic;
	 signal  berase_opcode :	std_logic_vector (7 downto 0);
	 signal  bp0_wire :	std_logic;
	 signal  bp1_wire :	std_logic;
	 signal  bp2_wire :	std_logic;
	 signal  bp3_wire :	std_logic;
	 signal  busy_wire :	std_logic;
	 signal  clkin_wire :	std_logic;
	 signal  clr_addmsb_wire :	std_logic;
	 signal  clr_endrbyte_wire :	std_logic;
	 signal  clr_read_wire :	std_logic;
	 signal  clr_read_wire2 :	std_logic;
	 signal  clr_rstat_wire :	std_logic;
	 signal  clr_write_wire :	std_logic;
	 signal  clr_write_wire2 :	std_logic;
	 signal  data0out_wire :	std_logic;
	 signal  data_valid_wire :	std_logic;
	 signal  datain_reg_wire_in :	std_logic_vector (7 downto 0);
	 signal  datain_wire :	std_logic_vector (3 downto 0);
	 signal  dataout_wire :	std_logic_vector (3 downto 0);
	 signal  derase_opcode :	std_logic_vector (7 downto 0);
	 signal  do_4baddr :	std_logic;
	 signal  do_bulk_erase :	std_logic;
	 signal  do_die_erase :	std_logic;
	 signal  do_ex4baddr :	std_logic;
	 signal  do_fast_read :	std_logic;
	 signal  do_fread_epcq :	std_logic;
	 signal  do_freadwrv_polling :	std_logic;
	 signal  do_memadd :	std_logic;
	 signal  do_polling :	std_logic;
	 signal  do_read :	std_logic;
	 signal  do_read_nonvolatile :	std_logic;
	 signal  do_read_rdid :	std_logic;
	 signal  do_read_sid :	std_logic;
	 signal  do_read_stat :	std_logic;
	 signal  do_read_volatile :	std_logic;
	 signal  do_sec_erase :	std_logic;
	 signal  do_sec_prot :	std_logic;
	 signal  do_secprot_wren :	std_logic;
	 signal  do_sprot_polling :	std_logic;
	 signal  do_sprot_rstat :	std_logic;
	 signal  do_wait_dummyclk :	std_logic;
	 signal  do_wren :	std_logic;
	 signal  do_write :	std_logic;
	 signal  do_write_polling :	std_logic;
	 signal  do_write_rstat :	std_logic;
	 signal  do_write_volatile :	std_logic;
	 signal  do_write_volatile_rstat :	std_logic;
	 signal  do_write_volatile_wren :	std_logic;
	 signal  do_write_wren :	std_logic;
	 signal  end1_cyc_gen_cntr_wire :	std_logic;
	 signal  end1_cyc_normal_in_wire :	std_logic;
	 signal  end1_cyc_reg_in_wire :	std_logic;
	 signal  end_add_cycle :	std_logic;
	 signal  end_add_cycle_mux_datab_wire :	std_logic;
	 signal  end_fast_read :	std_logic;
	 signal  end_one_cyc_pos :	std_logic;
	 signal  end_one_cycle :	std_logic;
	 signal  end_op_wire :	std_logic;
	 signal  end_operation :	std_logic;
	 signal  end_ophdly :	std_logic;
	 signal  end_pgwr_data :	std_logic;
	 signal  end_read :	std_logic;
	 signal  end_read_byte :	std_logic;
	 signal  end_wrstage :	std_logic;
	 signal  exb4addr_opcode :	std_logic_vector (7 downto 0);
	 signal  fast_read_opcode :	std_logic_vector (7 downto 0);
	 signal  fast_read_wire :	std_logic;
	 signal  freadwrv_sdoin :	std_logic;
	 signal  ill_write_wire :	std_logic;
	 signal  illegal_write_b4out_wire :	std_logic;
	 signal  illegal_write_prot :	std_logic;
	 signal  in_operation :	std_logic;
	 signal  load_opcode :	std_logic;
	 signal  mask_prot :	std_logic_vector (2 downto 0);
	 signal  mask_prot_add :	std_logic_vector (2 downto 0);
	 signal  mask_prot_check :	std_logic_vector (2 downto 0);
	 signal  mask_prot_comp_ntb :	std_logic_vector (2 downto 0);
	 signal  mask_prot_comp_tb :	std_logic_vector (2 downto 0);
	 signal  memadd_sdoin :	std_logic;
	 signal  ncs_reg_ena_wire :	std_logic;
	 signal  not_busy :	std_logic;
	 signal  oe_wire :	std_logic;
	 signal  pagewr_buf_not_empty :	std_logic_vector (0 downto 0);
	 signal  prot_wire :	std_logic_vector (7 downto 0);
	 signal  rden_wire :	std_logic;
	 signal  rdid_opcode :	std_logic_vector (7 downto 0);
	 signal  rdummyclk_opcode :	std_logic_vector (7 downto 0);
	 signal  read_data_reg_in_wire :	std_logic_vector (7 downto 0);
	 signal  read_opcode :	std_logic_vector (7 downto 0);
	 signal  read_rdid_wire :	std_logic;
	 signal  read_sid_wire :	std_logic;
	 signal  read_status_wire :	std_logic;
	 signal  read_wire :	std_logic;
	 signal  rflagstat_opcode :	std_logic_vector (7 downto 0);
	 signal  rnvdummyclk_opcode :	std_logic_vector (7 downto 0);
	 signal  rsid_opcode :	std_logic_vector (7 downto 0);
	 signal  rsid_sdoin :	std_logic;
	 signal  rstat_opcode :	std_logic_vector (7 downto 0);
	 signal  scein_wire :	std_logic;
	 signal  sdoin_wire :	std_logic;
	 signal  sec_protect_wire :	std_logic;
	 signal  secprot_opcode :	std_logic_vector (7 downto 0);
	 signal  secprot_sdoin :	std_logic;
	 signal  serase_opcode :	std_logic_vector (7 downto 0);
	 signal  shift_opcode :	std_logic;
	 signal  shift_opdata :	std_logic;
	 signal  shift_pgwr_data :	std_logic;
	 signal  st_busy_wire :	std_logic;
	 signal  stage2_wire :	std_logic;
	 signal  stage3_wire :	std_logic;
	 signal  stage4_wire :	std_logic;
	 signal  start_frpoll :	std_logic;
	 signal  start_poll :	std_logic;
	 signal  start_sppoll :	std_logic;
	 signal  start_wrpoll :	std_logic;
	 signal  to_sdoin_wire :	std_logic;
	 signal  wren_opcode :	std_logic_vector (7 downto 0);
	 signal  wren_wire :	std_logic;
	 signal  write_opcode :	std_logic_vector (7 downto 0);
	 signal  write_prot_true :	std_logic;
	 signal  write_prot_true2 :	std_logic;
	 signal  write_sdoin :	std_logic;
	 signal  write_wire :	std_logic;
	 signal  wrvolatile_opcode :	std_logic_vector (7 downto 0);
	 signal  wire_w_addr_range403w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_addr_range395w	:	std_logic_vector (22 downto 0);
	 signal  wire_w_addr_reg_overdie_range401w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_addr_reg_overdie_range391w	:	std_logic_vector (22 downto 0);
	 signal  wire_w_b4addr_opcode_range266w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_b4addr_opcode_range175w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_berase_opcode_range270w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_berase_opcode_range183w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_datain_range621w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_datain_range616w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_dataout_wire_range445w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_derase_opcode_range272w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_derase_opcode_range188w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_exb4addr_opcode_range264w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_exb4addr_opcode_range170w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_fast_read_opcode_range288w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_fast_read_opcode_range228w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_mask_prot_range568w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_mask_prot_range571w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_mask_prot_range573w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_mask_prot_add_range576w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_mask_prot_add_range583w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_mask_prot_add_range588w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_mask_prot_check_range585w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_mask_prot_check_range590w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_mask_prot_comp_ntb_range591w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_mask_prot_comp_ntb_range596w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_mask_prot_comp_tb_range593w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_mask_prot_comp_tb_range598w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_pagewr_buf_not_empty_range68w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_prot_wire_range551w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_prot_wire_range553w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_prot_wire_range556w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_rdid_opcode_range294w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_rdid_opcode_range239w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_rdummyclk_opcode_range286w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_rdummyclk_opcode_range221w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_read_opcode_range290w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_read_opcode_range231w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_rflagstat_opcode_range276w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_rflagstat_opcode_range198w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_rnvdummyclk_opcode_range282w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_rnvdummyclk_opcode_range211w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_rsid_opcode_range296w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_rsid_opcode_range242w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_rstat_opcode_range278w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_rstat_opcode_range202w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_secprot_opcode_range292w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_secprot_opcode_range234w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_serase_opcode_range274w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_serase_opcode_range193w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_wren_opcode_range268w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_wren_opcode_range180w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_write_opcode_range280w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_write_opcode_range206w	:	std_logic_vector (6 downto 0);
	 signal  wire_w_wrvolatile_opcode_range284w	:	std_logic_vector (0 downto 0);
	 signal  wire_w_wrvolatile_opcode_range214w	:	std_logic_vector (6 downto 0);
	 component  a_graycounter
	 generic 
	 (
		pvalue	:	natural := 0;
		width	:	natural := 8;
		lpm_type	:	string := "a_graycounter"
	 );
	 port
	 ( 
		aclr	:	in std_logic := '0';
		clk_en	:	in std_logic := '1';
		clock	:	in std_logic;
		cnt_en	:	in std_logic := '1';
		q	:	out std_logic_vector(width-1 downto 0);
		qbin	:	out std_logic_vector(width-1 downto 0);
		sclr	:	in std_logic := '0';
		updown	:	in std_logic := '1'
	 ); 
	 end component;
	 component  cycloneii_asmiblock
	 port
	 ( 
		data0out	:	out std_logic;
		dclkin	:	in std_logic;
		oe	:	in std_logic := '1';
		scein	:	in std_logic;
		sdoin	:	in std_logic
	 ); 
	 end component;
 begin

	wire_w_lg_w_lg_w655w656w657w(0) <= wire_w_lg_w655w656w(0) and end_operation;
	wire_w_lg_w655w656w(0) <= wire_w655w(0) and wire_w_lg_do_ex4baddr646w(0);
	wire_w287w(0) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode223w224w225w226w(0) and wire_w_rdummyclk_opcode_range286w(0);
	loop0 : for i in 0 to 6 generate 
		wire_w227w(i) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode223w224w225w226w(0) and wire_w_rdummyclk_opcode_range221w(i);
	end generate loop0;
	wire_w285w(0) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode216w217w218w219w(0) and wire_w_wrvolatile_opcode_range284w(0);
	loop1 : for i in 0 to 6 generate 
		wire_w220w(i) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode216w217w218w219w(0) and wire_w_wrvolatile_opcode_range214w(i);
	end generate loop1;
	wire_w655w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_write651w652w653w654w(0) and wire_w_lg_do_4baddr647w(0);
	wire_w477w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_read407w474w475w476w(0) and end_read_byte;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode184w185w186w271w(0) <= wire_w_lg_w_lg_w_lg_load_opcode184w185w186w(0) and wire_w_berase_opcode_range270w(0);
	loop2 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode184w185w186w187w(i) <= wire_w_lg_w_lg_w_lg_load_opcode184w185w186w(0) and wire_w_berase_opcode_range183w(i);
	end generate loop2;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode189w190w191w273w(0) <= wire_w_lg_w_lg_w_lg_load_opcode189w190w191w(0) and wire_w_derase_opcode_range272w(0);
	loop3 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode189w190w191w192w(i) <= wire_w_lg_w_lg_w_lg_load_opcode189w190w191w(0) and wire_w_derase_opcode_range188w(i);
	end generate loop3;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode223w224w225w226w(0) <= wire_w_lg_w_lg_w_lg_load_opcode223w224w225w(0) and wire_w_lg_do_read_stat52w(0);
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode194w195w196w275w(0) <= wire_w_lg_w_lg_w_lg_load_opcode194w195w196w(0) and wire_w_serase_opcode_range274w(0);
	loop4 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode194w195w196w197w(i) <= wire_w_lg_w_lg_w_lg_load_opcode194w195w196w(0) and wire_w_serase_opcode_range193w(i);
	end generate loop4;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode235w236w237w293w(0) <= wire_w_lg_w_lg_w_lg_load_opcode235w236w237w(0) and wire_w_secprot_opcode_range292w(0);
	loop5 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode235w236w237w238w(i) <= wire_w_lg_w_lg_w_lg_load_opcode235w236w237w(0) and wire_w_secprot_opcode_range234w(i);
	end generate loop5;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode216w217w218w219w(0) <= wire_w_lg_w_lg_w_lg_load_opcode216w217w218w(0) and wire_w_lg_do_read_stat52w(0);
	wire_w_lg_w_lg_w_lg_w_lg_do_read359w360w361w362w(0) <= wire_w_lg_w_lg_w_lg_do_read359w360w361w(0) and end_one_cycle;
	wire_w_lg_w_lg_w_lg_w_lg_do_write651w652w653w654w(0) <= wire_w_lg_w_lg_w_lg_do_write651w652w653w(0) and wire_w_lg_do_die_erase648w(0);
	wire_w_lg_w_lg_w_lg_w530w641w642w658w(0) <= wire_w_lg_w_lg_w530w641w642w(0) and end_operation;
	wire_w_lg_w_lg_w_lg_w_lg_do_read407w474w475w476w(0) <= wire_w_lg_w_lg_w_lg_do_read407w474w475w(0) and end_one_cyc_pos;
	wire_w_lg_w_lg_w_lg_w_lg_do_sec_erase54w416w417w418w(0) <= wire_w_lg_w_lg_w_lg_do_sec_erase54w416w417w(0) and end_operation;
	wire_w_lg_w_lg_w_lg_do_write628w629w630w(0) <= wire_w_lg_w_lg_do_write628w629w(0) and stage4_wire;
	wire_w_lg_w_lg_w_lg_load_opcode184w185w186w(0) <= wire_w_lg_w_lg_load_opcode184w185w(0) and wire_w_lg_do_read_stat52w(0);
	wire_w_lg_w_lg_w_lg_load_opcode189w190w191w(0) <= wire_w_lg_w_lg_load_opcode189w190w(0) and wire_w_lg_do_read_stat52w(0);
	wire_w_lg_w_lg_w_lg_load_opcode199w204w279w(0) <= wire_w_lg_w_lg_load_opcode199w204w(0) and wire_w_rstat_opcode_range278w(0);
	loop6 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_w_lg_load_opcode199w204w205w(i) <= wire_w_lg_w_lg_load_opcode199w204w(0) and wire_w_rstat_opcode_range202w(i);
	end generate loop6;
	wire_w_lg_w_lg_w_lg_load_opcode199w200w277w(0) <= wire_w_lg_w_lg_load_opcode199w200w(0) and wire_w_rflagstat_opcode_range276w(0);
	loop7 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_w_lg_load_opcode199w200w201w(i) <= wire_w_lg_w_lg_load_opcode199w200w(0) and wire_w_rflagstat_opcode_range198w(i);
	end generate loop7;
	wire_w_lg_w_lg_w_lg_load_opcode223w224w225w(0) <= wire_w_lg_w_lg_load_opcode223w224w(0) and wire_w_lg_do_wren53w(0);
	wire_w_lg_w_lg_w_lg_load_opcode194w195w196w(0) <= wire_w_lg_w_lg_load_opcode194w195w(0) and wire_w_lg_do_read_stat52w(0);
	wire_w_lg_w_lg_w_lg_load_opcode235w236w237w(0) <= wire_w_lg_w_lg_load_opcode235w236w(0) and wire_w_lg_do_read_stat52w(0);
	wire_w_lg_w_lg_w_lg_load_opcode216w217w218w(0) <= wire_w_lg_w_lg_load_opcode216w217w(0) and wire_w_lg_do_wren53w(0);
	wire_w_lg_w_lg_w_lg_bp2_wire547w548w549w(0) <= wire_w_lg_w_lg_bp2_wire547w548w(0) and wire_w_lg_bp0_wire545w(0);
	wire_w_lg_w_lg_w_lg_bp2_wire547w548w552w(0) <= wire_w_lg_w_lg_bp2_wire547w548w(0) and bp0_wire;
	wire_w_lg_w_lg_w_lg_bp2_wire547w554w555w(0) <= wire_w_lg_w_lg_bp2_wire547w554w(0) and wire_w_lg_bp0_wire545w(0);
	wire_w_lg_w_lg_w_lg_bp2_wire547w554w557w(0) <= wire_w_lg_w_lg_bp2_wire547w554w(0) and bp0_wire;
	wire_w_lg_w_lg_w_lg_do_read359w360w361w(0) <= wire_w_lg_w_lg_do_read359w360w(0) and wire_w_lg_w_lg_do_write63w357w(0);
	wire_w_lg_w_lg_w_lg_do_read359w360w419w(0) <= wire_w_lg_w_lg_do_read359w360w(0) and clr_write_wire2;
	wire_w_lg_w_lg_w_lg_do_write651w652w653w(0) <= wire_w_lg_w_lg_do_write651w652w(0) and wire_w_lg_do_bulk_erase649w(0);
	wire_w_lg_w_lg_w530w641w642w(0) <= wire_w_lg_w530w641w(0) and wire_wrstage_cntr_w_lg_w_q_range522w523w(0);
	wire_w_lg_w_lg_w_lg_do_read407w474w475w(0) <= wire_w_lg_w_lg_do_read407w474w(0) and wire_stage_cntr_w_lg_w_q_range102w107w(0);
	wire_w_lg_w_lg_w_lg_do_sec_erase54w416w417w(0) <= wire_w_lg_w_lg_do_sec_erase54w416w(0) and wire_w_lg_do_read_stat52w(0);
	wire_w_lg_w_lg_bp2_wire559w560w(0) <= wire_w_lg_bp2_wire559w(0) and wire_w_lg_bp0_wire545w(0);
	wire_w_lg_w_lg_bp2_wire559w562w(0) <= wire_w_lg_bp2_wire559w(0) and bp0_wire;
	wire_w_lg_w_lg_bp2_wire564w565w(0) <= wire_w_lg_bp2_wire564w(0) and wire_w_lg_bp0_wire545w(0);
	wire_w_lg_w_lg_bp2_wire564w567w(0) <= wire_w_lg_bp2_wire564w(0) and bp0_wire;
	wire_w_lg_w_lg_do_4baddr176w177w(0) <= wire_w_lg_do_4baddr176w(0) and wire_w_lg_do_wren53w(0);
	wire_w_lg_w_lg_do_ex4baddr171w172w(0) <= wire_w_lg_do_ex4baddr171w(0) and wire_w_lg_do_wren53w(0);
	wire_w_lg_w_lg_do_polling500w501w(0) <= wire_w_lg_do_polling500w(0) and stage3_dly_reg;
	wire_w_lg_w_lg_do_read_stat123w124w(0) <= wire_w_lg_do_read_stat123w(0) and wire_w_lg_w_lg_w119w120w121w(0);
	wire_w_lg_w_lg_do_write207w208w(0) <= wire_w_lg_do_write207w(0) and wire_w_lg_do_wren53w(0);
	wire_w_lg_w_lg_do_write628w629w(0) <= wire_w_lg_do_write628w(0) and wire_w_lg_do_write_rstat627w(0);
	wire_w_lg_w_lg_do_write63w338w(0) <= wire_w_lg_do_write63w(0) and end_pgwr_data;
	wire_w_lg_w_lg_load_opcode178w267w(0) <= wire_w_lg_load_opcode178w(0) and wire_w_b4addr_opcode_range266w(0);
	loop8 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_load_opcode178w179w(i) <= wire_w_lg_load_opcode178w(0) and wire_w_b4addr_opcode_range175w(i);
	end generate loop8;
	wire_w_lg_w_lg_load_opcode173w265w(0) <= wire_w_lg_load_opcode173w(0) and wire_w_exb4addr_opcode_range264w(0);
	loop9 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_load_opcode173w174w(i) <= wire_w_lg_load_opcode173w(0) and wire_w_exb4addr_opcode_range170w(i);
	end generate loop9;
	wire_w_lg_w_lg_load_opcode209w281w(0) <= wire_w_lg_load_opcode209w(0) and wire_w_write_opcode_range280w(0);
	loop10 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_load_opcode209w210w(i) <= wire_w_lg_load_opcode209w(0) and wire_w_write_opcode_range206w(i);
	end generate loop10;
	wire_w_lg_w_lg_load_opcode184w185w(0) <= wire_w_lg_load_opcode184w(0) and wire_w_lg_do_wren53w(0);
	wire_w_lg_w_lg_load_opcode189w190w(0) <= wire_w_lg_load_opcode189w(0) and wire_w_lg_do_wren53w(0);
	wire_w_lg_w_lg_load_opcode229w289w(0) <= wire_w_lg_load_opcode229w(0) and wire_w_fast_read_opcode_range288w(0);
	loop11 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_load_opcode229w230w(i) <= wire_w_lg_load_opcode229w(0) and wire_w_fast_read_opcode_range228w(i);
	end generate loop11;
	wire_w_lg_w_lg_load_opcode232w291w(0) <= wire_w_lg_load_opcode232w(0) and wire_w_read_opcode_range290w(0);
	loop12 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_load_opcode232w233w(i) <= wire_w_lg_load_opcode232w(0) and wire_w_read_opcode_range231w(i);
	end generate loop12;
	wire_w_lg_w_lg_load_opcode212w283w(0) <= wire_w_lg_load_opcode212w(0) and wire_w_rnvdummyclk_opcode_range282w(0);
	loop13 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_load_opcode212w213w(i) <= wire_w_lg_load_opcode212w(0) and wire_w_rnvdummyclk_opcode_range211w(i);
	end generate loop13;
	wire_w_lg_w_lg_load_opcode240w295w(0) <= wire_w_lg_load_opcode240w(0) and wire_w_rdid_opcode_range294w(0);
	loop14 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_load_opcode240w241w(i) <= wire_w_lg_load_opcode240w(0) and wire_w_rdid_opcode_range239w(i);
	end generate loop14;
	wire_w_lg_w_lg_load_opcode243w297w(0) <= wire_w_lg_load_opcode243w(0) and wire_w_rsid_opcode_range296w(0);
	loop15 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_load_opcode243w244w(i) <= wire_w_lg_load_opcode243w(0) and wire_w_rsid_opcode_range242w(i);
	end generate loop15;
	wire_w_lg_w_lg_load_opcode199w204w(0) <= wire_w_lg_load_opcode199w(0) and wire_w_lg_do_polling203w(0);
	wire_w_lg_w_lg_load_opcode199w200w(0) <= wire_w_lg_load_opcode199w(0) and do_polling;
	wire_w_lg_w_lg_load_opcode223w224w(0) <= wire_w_lg_load_opcode223w(0) and wire_w_lg_do_write_volatile222w(0);
	wire_w_lg_w_lg_load_opcode194w195w(0) <= wire_w_lg_load_opcode194w(0) and wire_w_lg_do_wren53w(0);
	wire_w_lg_w_lg_load_opcode235w236w(0) <= wire_w_lg_load_opcode235w(0) and wire_w_lg_do_wren53w(0);
	wire_w_lg_w_lg_load_opcode181w269w(0) <= wire_w_lg_load_opcode181w(0) and wire_w_wren_opcode_range268w(0);
	loop16 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_load_opcode181w182w(i) <= wire_w_lg_load_opcode181w(0) and wire_w_wren_opcode_range180w(i);
	end generate loop16;
	wire_w_lg_w_lg_load_opcode216w217w(0) <= wire_w_lg_load_opcode216w(0) and wire_w_lg_do_read_volatile215w(0);
	wire_w_lg_w_lg_stage3_wire45w46w(0) <= wire_w_lg_stage3_wire45w(0) and do_wait_dummyclk;
	wire_w_lg_w_lg_start_poll345w346w(0) <= wire_w_lg_start_poll345w(0) and do_polling;
	wire_w_lg_w_lg_bp2_wire547w548w(0) <= wire_w_lg_bp2_wire547w(0) and wire_w_lg_bp1_wire546w(0);
	wire_w_lg_w_lg_bp2_wire547w554w(0) <= wire_w_lg_bp2_wire547w(0) and bp1_wire;
	wire_w_lg_w_lg_do_read359w360w(0) <= wire_w_lg_do_read359w(0) and wire_w_lg_do_fast_read358w(0);
	wire_w_lg_w_lg_do_write651w652w(0) <= wire_w_lg_do_write651w(0) and wire_w_lg_do_sec_erase650w(0);
	wire_w_lg_w_lg_w517w518w519w(0) <= wire_w_lg_w517w518w(0) and end_wrstage;
	wire_w_lg_w530w641w(0) <= wire_w530w(0) and wire_wrstage_cntr_w_q_range524w(0);
	wire_w_lg_w_lg_w_lg_w_lg_do_write72w116w117w516w(0) <= wire_w_lg_w_lg_w_lg_do_write72w116w117w(0) and wire_w_lg_write_prot_true515w(0);
	wire_w_lg_w_lg_w_lg_w_lg_do_write72w116w117w130w(0) <= wire_w_lg_w_lg_w_lg_do_write72w116w117w(0) and write_prot_true;
	wire_w_lg_w_lg_w_lg_do_write72w73w408w(0) <= wire_w_lg_w_lg_do_write72w73w(0) and do_memadd;
	wire_w_lg_w_lg_do_read407w474w(0) <= wire_w_lg_do_read407w(0) and wire_stage_cntr_w_q_range103w(0);
	wire_w_lg_w_lg_do_read_rdid125w126w(0) <= wire_w_lg_do_read_rdid125w(0) and end_op_wire;
	wire_w_lg_w_lg_do_sec_erase54w416w(0) <= wire_w_lg_do_sec_erase54w(0) and wire_w_lg_do_wren53w(0);
	wire_w_lg_w_lg_end_operation502w503w(0) <= wire_w_lg_end_operation502w(0) and do_read_stat;
	wire_w_lg_w_lg_rden_wire412w413w(0) <= wire_w_lg_rden_wire412w(0) and not_busy;
	wire_w_lg_addr_overdie402w(0) <= addr_overdie and wire_w_addr_reg_overdie_range401w(0);
	loop17 : for i in 0 to 22 generate 
		wire_w_lg_addr_overdie392w(i) <= addr_overdie and wire_w_addr_reg_overdie_range391w(i);
	end generate loop17;
	wire_w_lg_bp2_wire559w(0) <= bp2_wire and wire_w_lg_bp1_wire546w(0);
	wire_w_lg_bp2_wire564w(0) <= bp2_wire and bp1_wire;
	wire_w_lg_do_4baddr176w(0) <= do_4baddr and wire_w_lg_do_read_stat52w(0);
	wire_w_lg_do_bulk_erase339w(0) <= do_bulk_erase and wire_w_lg_do_read_stat52w(0);
	wire_w_lg_do_ex4baddr171w(0) <= do_ex4baddr and wire_w_lg_do_read_stat52w(0);
	wire_w_lg_do_polling500w(0) <= do_polling and end_one_cyc_pos;
	wire_w_lg_do_read_nonvolatile325w(0) <= do_read_nonvolatile and wire_addbyte_cntr_w_q_range158w(0);
	wire_w_lg_do_read_stat123w(0) <= do_read_stat and wire_w_lg_start_poll122w(0);
	wire_w_lg_do_write207w(0) <= do_write and wire_w_lg_do_read_stat52w(0);
	wire_w_lg_do_write628w(0) <= do_write and wire_w_lg_do_wren53w(0);
	wire_w_lg_do_write70w(0) <= do_write and wire_w_lg_w_pagewr_buf_not_empty_range68w69w(0);
	wire_w_lg_do_write63w(0) <= do_write and shift_pgwr_data;
	wire_w_lg_load_opcode178w(0) <= load_opcode and wire_w_lg_w_lg_do_4baddr176w177w(0);
	wire_w_lg_load_opcode173w(0) <= load_opcode and wire_w_lg_w_lg_do_ex4baddr171w172w(0);
	wire_w_lg_load_opcode209w(0) <= load_opcode and wire_w_lg_w_lg_do_write207w208w(0);
	wire_w_lg_load_opcode184w(0) <= load_opcode and do_bulk_erase;
	wire_w_lg_load_opcode189w(0) <= load_opcode and do_die_erase;
	wire_w_lg_load_opcode229w(0) <= load_opcode and do_fast_read;
	wire_w_lg_load_opcode232w(0) <= load_opcode and do_read;
	wire_w_lg_load_opcode212w(0) <= load_opcode and do_read_nonvolatile;
	wire_w_lg_load_opcode240w(0) <= load_opcode and do_read_rdid;
	wire_w_lg_load_opcode243w(0) <= load_opcode and do_read_sid;
	wire_w_lg_load_opcode199w(0) <= load_opcode and do_read_stat;
	wire_w_lg_load_opcode223w(0) <= load_opcode and do_read_volatile;
	wire_w_lg_load_opcode194w(0) <= load_opcode and do_sec_erase;
	wire_w_lg_load_opcode235w(0) <= load_opcode and do_sec_prot;
	wire_w_lg_load_opcode181w(0) <= load_opcode and do_wren;
	wire_w_lg_load_opcode216w(0) <= load_opcode and do_write_volatile;
	wire_w_lg_not_busy404w(0) <= not_busy and wire_w_addr_range403w(0);
	loop18 : for i in 0 to 22 generate 
		wire_w_lg_not_busy396w(i) <= not_busy and wire_w_addr_range395w(i);
	end generate loop18;
	wire_w_lg_not_busy622w(0) <= not_busy and wire_w_datain_range621w(0);
	loop19 : for i in 0 to 6 generate 
		wire_w_lg_not_busy617w(i) <= not_busy and wire_w_datain_range616w(i);
	end generate loop19;
	loop20 : for i in 0 to 6 generate 
		wire_w_lg_shift_opcode169w(i) <= shift_opcode and wire_asmi_opcode_reg_w_q_range168w(i);
	end generate loop20;
	wire_w_lg_stage3_wire410w(0) <= stage3_wire and wire_w_lg_w_lg_w_lg_w_lg_do_write72w73w408w409w(0);
	wire_w_lg_stage3_wire441w(0) <= stage3_wire and wire_w_lg_w_lg_w_lg_do_read_stat438w439w440w(0);
	wire_w_lg_stage3_wire55w(0) <= stage3_wire and wire_w_lg_do_sec_erase54w(0);
	wire_w_lg_stage3_wire45w(0) <= stage3_wire and do_fast_read;
	loop21 : for i in 0 to 22 generate 
		wire_w_lg_stage3_wire394w(i) <= stage3_wire and wire_addr_reg_w_q_range393w(i);
	end generate loop21;
	wire_w_lg_stage4_wire443w(0) <= stage4_wire and wire_w_lg_w_lg_do_read407w442w(0);
	wire_w_lg_stage4_wire411w(0) <= stage4_wire and addr_overdie;
	loop22 : for i in 0 to 6 generate 
		wire_w_lg_stage4_wire615w(i) <= stage4_wire and wire_datain_reg_w_q_range614w(i);
	end generate loop22;
	wire_w_lg_start_poll345w(0) <= start_poll and do_read_stat;
	wire_w_lg_wren_wire631w(0) <= wren_wire and not_busy;
	wire_w_lg_w_mask_prot_range568w575w(0) <= wire_w_mask_prot_range568w(0) and wire_addr_reg_w_q_range574w(0);
	wire_w_lg_w_mask_prot_range571w582w(0) <= wire_w_mask_prot_range571w(0) and wire_addr_reg_w_q_range581w(0);
	wire_w_lg_w_mask_prot_range573w587w(0) <= wire_w_mask_prot_range573w(0) and wire_addr_reg_w_q_range586w(0);
	wire_w_lg_w_lg_do_write63w357w(0) <= not wire_w_lg_do_write63w(0);
	wire_w_lg_w_lg_w119w120w121w(0) <= not wire_w_lg_w119w120w(0);
	wire_w_lg_addr_overdie490w(0) <= not addr_overdie;
	wire_w_lg_bp0_wire545w(0) <= not bp0_wire;
	wire_w_lg_bp1_wire546w(0) <= not bp1_wire;
	wire_w_lg_bp2_wire547w(0) <= not bp2_wire;
	wire_w_lg_busy_wire1w(0) <= not busy_wire;
	wire_w_lg_clkin_wire101w(0) <= not clkin_wire;
	wire_w_lg_do_4baddr647w(0) <= not do_4baddr;
	wire_w_lg_do_bulk_erase649w(0) <= not do_bulk_erase;
	wire_w_lg_do_die_erase648w(0) <= not do_die_erase;
	wire_w_lg_do_ex4baddr646w(0) <= not do_ex4baddr;
	wire_w_lg_do_fast_read358w(0) <= not do_fast_read;
	wire_w_lg_do_memadd425w(0) <= not do_memadd;
	wire_w_lg_do_polling203w(0) <= not do_polling;
	wire_w_lg_do_read359w(0) <= not do_read;
	wire_w_lg_do_read_rdid51w(0) <= not do_read_rdid;
	wire_w_lg_do_read_stat52w(0) <= not do_read_stat;
	wire_w_lg_do_read_volatile215w(0) <= not do_read_volatile;
	wire_w_lg_do_sec_erase650w(0) <= not do_sec_erase;
	wire_w_lg_do_wren53w(0) <= not do_wren;
	wire_w_lg_do_write651w(0) <= not do_write;
	wire_w_lg_do_write_rstat627w(0) <= not do_write_rstat;
	wire_w_lg_do_write_volatile222w(0) <= not do_write_volatile;
	wire_w_lg_end_add_cycle83w(0) <= not end_add_cycle;
	wire_w_lg_end_fast_read77w(0) <= not end_fast_read;
	wire_w_lg_end_ophdly39w(0) <= not end_ophdly;
	wire_w_lg_end_pgwr_data62w(0) <= not end_pgwr_data;
	wire_w_lg_end_read80w(0) <= not end_read;
	wire_w_lg_rden_wire492w(0) <= not rden_wire;
	wire_w_lg_read_rdid_wire9w(0) <= not read_rdid_wire;
	wire_w_lg_read_sid_wire8w(0) <= not read_sid_wire;
	wire_w_lg_sec_protect_wire7w(0) <= not sec_protect_wire;
	wire_w_lg_st_busy_wire127w(0) <= not st_busy_wire;
	wire_w_lg_start_poll122w(0) <= not start_poll;
	wire_w_lg_write_prot_true515w(0) <= not write_prot_true;
	wire_w_lg_write_wire17w(0) <= not write_wire;
	wire_w_lg_w_pagewr_buf_not_empty_range68w69w(0) <= not wire_w_pagewr_buf_not_empty_range68w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w530w641w642w658w659w(0) <= wire_w_lg_w_lg_w_lg_w530w641w642w658w(0) or write_prot_true;
	wire_w_lg_w_lg_w_lg_load_opcode243w297w298w(0) <= wire_w_lg_w_lg_load_opcode243w297w(0) or wire_w_lg_w_lg_load_opcode240w295w(0);
	loop23 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_w_lg_load_opcode243w244w245w(i) <= wire_w_lg_w_lg_load_opcode243w244w(i) or wire_w_lg_w_lg_load_opcode240w241w(i);
	end generate loop23;
	wire_w517w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_write72w116w117w516w(0) or do_4baddr;
	wire_w_lg_w_lg_w_lg_w_lg_do_write72w73w408w409w(0) <= wire_w_lg_w_lg_w_lg_do_write72w73w408w(0) or wire_w_lg_do_read407w(0);
	wire_w_lg_w_lg_w_lg_end_operation502w503w504w(0) <= wire_w_lg_w_lg_end_operation502w503w(0) or clr_rstat_wire;
	wire_w_lg_w_lg_w_lg_rden_wire412w413w414w(0) <= wire_w_lg_w_lg_rden_wire412w413w(0) or wire_w_lg_stage4_wire411w(0);
	wire_w_lg_w_lg_not_busy404w405w(0) <= wire_w_lg_not_busy404w(0) or wire_w_lg_addr_overdie402w(0);
	loop24 : for i in 0 to 22 generate 
		wire_w_lg_w_lg_not_busy396w397w(i) <= wire_w_lg_not_busy396w(i) or wire_w_lg_stage3_wire394w(i);
	end generate loop24;
	loop25 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_not_busy617w618w(i) <= wire_w_lg_not_busy617w(i) or wire_w_lg_stage4_wire615w(i);
	end generate loop25;
	wire_w_lg_w_lg_stage4_wire443w444w(0) <= wire_w_lg_stage4_wire443w(0) or wire_w_lg_stage3_wire441w(0);
	wire_w_lg_w_lg_wren_wire631w632w(0) <= wire_w_lg_wren_wire631w(0) or wire_w_lg_w_lg_w_lg_do_write628w629w630w(0);
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode243w297w298w299w(0) <= wire_w_lg_w_lg_w_lg_load_opcode243w297w298w(0) or wire_w_lg_w_lg_w_lg_w_lg_load_opcode235w236w237w293w(0);
	loop26 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode243w244w245w246w(i) <= wire_w_lg_w_lg_w_lg_load_opcode243w244w245w(i) or wire_w_lg_w_lg_w_lg_w_lg_load_opcode235w236w237w238w(i);
	end generate loop26;
	wire_w_lg_w517w518w(0) <= wire_w517w(0) or do_ex4baddr;
	wire_w_lg_w_lg_w_lg_w_lg_rden_wire412w413w414w415w(0) <= wire_w_lg_w_lg_w_lg_rden_wire412w413w414w(0) or wire_w_lg_stage3_wire410w(0);
	loop27 : for i in 0 to 22 generate 
		wire_w_lg_w_lg_w_lg_not_busy396w397w398w(i) <= wire_w_lg_w_lg_not_busy396w397w(i) or wire_w_lg_addr_overdie392w(i);
	end generate loop27;
	wire_w300w(0) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode243w297w298w299w(0) or wire_w_lg_w_lg_load_opcode232w291w(0);
	loop28 : for i in 0 to 6 generate 
		wire_w247w(i) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode243w244w245w246w(i) or wire_w_lg_w_lg_load_opcode232w233w(i);
	end generate loop28;
	wire_w_lg_w300w301w(0) <= wire_w300w(0) or wire_w_lg_w_lg_load_opcode229w289w(0);
	loop29 : for i in 0 to 6 generate 
		wire_w_lg_w247w248w(i) <= wire_w247w(i) or wire_w_lg_w_lg_load_opcode229w230w(i);
	end generate loop29;
	wire_w_lg_w_lg_w300w301w302w(0) <= wire_w_lg_w300w301w(0) or wire_w287w(0);
	loop30 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_w247w248w249w(i) <= wire_w_lg_w247w248w(i) or wire_w227w(i);
	end generate loop30;
	wire_w_lg_w_lg_w_lg_w300w301w302w303w(0) <= wire_w_lg_w_lg_w300w301w302w(0) or wire_w285w(0);
	loop31 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_w_lg_w247w248w249w250w(i) <= wire_w_lg_w_lg_w247w248w249w(i) or wire_w220w(i);
	end generate loop31;
	wire_w_lg_w_lg_w_lg_w_lg_w300w301w302w303w304w(0) <= wire_w_lg_w_lg_w_lg_w300w301w302w303w(0) or wire_w_lg_w_lg_load_opcode212w283w(0);
	loop32 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_w_lg_w_lg_w247w248w249w250w251w(i) <= wire_w_lg_w_lg_w_lg_w247w248w249w250w(i) or wire_w_lg_w_lg_load_opcode212w213w(i);
	end generate loop32;
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w300w301w302w303w304w305w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w300w301w302w303w304w(0) or wire_w_lg_w_lg_load_opcode209w281w(0);
	loop33 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_w_lg_w_lg_w_lg_w247w248w249w250w251w252w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w247w248w249w250w251w(i) or wire_w_lg_w_lg_load_opcode209w210w(i);
	end generate loop33;
	wire_w306w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w300w301w302w303w304w305w(0) or wire_w_lg_w_lg_w_lg_load_opcode199w204w279w(0);
	loop34 : for i in 0 to 6 generate 
		wire_w253w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w247w248w249w250w251w252w(i) or wire_w_lg_w_lg_w_lg_load_opcode199w204w205w(i);
	end generate loop34;
	wire_w_lg_w306w307w(0) <= wire_w306w(0) or wire_w_lg_w_lg_w_lg_load_opcode199w200w277w(0);
	loop35 : for i in 0 to 6 generate 
		wire_w_lg_w253w254w(i) <= wire_w253w(i) or wire_w_lg_w_lg_w_lg_load_opcode199w200w201w(i);
	end generate loop35;
	wire_w_lg_w_lg_w306w307w308w(0) <= wire_w_lg_w306w307w(0) or wire_w_lg_w_lg_w_lg_w_lg_load_opcode194w195w196w275w(0);
	loop36 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_w253w254w255w(i) <= wire_w_lg_w253w254w(i) or wire_w_lg_w_lg_w_lg_w_lg_load_opcode194w195w196w197w(i);
	end generate loop36;
	wire_w_lg_w_lg_w_lg_w306w307w308w309w(0) <= wire_w_lg_w_lg_w306w307w308w(0) or wire_w_lg_w_lg_w_lg_w_lg_load_opcode189w190w191w273w(0);
	loop37 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_w_lg_w253w254w255w256w(i) <= wire_w_lg_w_lg_w253w254w255w(i) or wire_w_lg_w_lg_w_lg_w_lg_load_opcode189w190w191w192w(i);
	end generate loop37;
	wire_w_lg_w_lg_w_lg_w_lg_w306w307w308w309w310w(0) <= wire_w_lg_w_lg_w_lg_w306w307w308w309w(0) or wire_w_lg_w_lg_w_lg_w_lg_load_opcode184w185w186w271w(0);
	loop38 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_w_lg_w_lg_w253w254w255w256w257w(i) <= wire_w_lg_w_lg_w_lg_w253w254w255w256w(i) or wire_w_lg_w_lg_w_lg_w_lg_load_opcode184w185w186w187w(i);
	end generate loop38;
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w306w307w308w309w310w311w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w306w307w308w309w310w(0) or wire_w_lg_w_lg_load_opcode181w269w(0);
	loop39 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_w_lg_w_lg_w_lg_w253w254w255w256w257w258w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w253w254w255w256w257w(i) or wire_w_lg_w_lg_load_opcode181w182w(i);
	end generate loop39;
	wire_w312w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w306w307w308w309w310w311w(0) or wire_w_lg_w_lg_load_opcode178w267w(0);
	loop40 : for i in 0 to 6 generate 
		wire_w259w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w253w254w255w256w257w258w(i) or wire_w_lg_w_lg_load_opcode178w179w(i);
	end generate loop40;
	wire_w_lg_w312w313w(0) <= wire_w312w(0) or wire_w_lg_w_lg_load_opcode173w265w(0);
	loop41 : for i in 0 to 6 generate 
		wire_w_lg_w259w260w(i) <= wire_w259w(i) or wire_w_lg_w_lg_load_opcode173w174w(i);
	end generate loop41;
	loop42 : for i in 0 to 6 generate 
		wire_w_lg_w_lg_w259w260w261w(i) <= wire_w_lg_w259w260w(i) or wire_w_lg_shift_opcode169w(i);
	end generate loop42;
	wire_w_lg_w_lg_w151w152w153w(0) <= wire_w_lg_w151w152w(0) or do_read_nonvolatile;
	wire_w_lg_w151w152w(0) <= wire_w151w(0) or do_fast_read;
	wire_w_lg_w119w120w(0) <= wire_w119w(0) or do_ex4baddr;
	wire_w151w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_read_sid147w148w149w150w(0) or do_read;
	wire_w530w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_write72w116w117w529w(0) or do_ex4baddr;
	wire_w119w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_write72w116w117w118w(0) or do_4baddr;
	wire_w_lg_w_lg_w_lg_w_lg_do_read407w428w429w430w(0) <= wire_w_lg_w_lg_w_lg_do_read407w428w429w(0) or do_die_erase;
	wire_w_lg_w_lg_w_lg_w_lg_do_read_sid147w148w149w150w(0) <= wire_w_lg_w_lg_w_lg_do_read_sid147w148w149w(0) or do_read_rdid;
	wire_w_lg_w_lg_w_lg_w_lg_do_write72w116w117w529w(0) <= wire_w_lg_w_lg_w_lg_do_write72w116w117w(0) or do_4baddr;
	wire_w_lg_w_lg_w_lg_w_lg_do_write72w116w117w118w(0) <= wire_w_lg_w_lg_w_lg_do_write72w116w117w(0) or do_fread_epcq;
	wire_w_lg_w_lg_w_lg_bp3_wire539w540w541w(0) <= wire_w_lg_w_lg_bp3_wire539w540w(0) or bp0_wire;
	wire_w_lg_w_lg_w_lg_do_read407w428w429w(0) <= wire_w_lg_w_lg_do_read407w428w(0) or do_sec_erase;
	wire_w_lg_w_lg_w_lg_do_read_sid147w148w149w(0) <= wire_w_lg_w_lg_do_read_sid147w148w(0) or do_die_erase;
	wire_w_lg_w_lg_w_lg_do_read_stat438w439w440w(0) <= wire_w_lg_w_lg_do_read_stat438w439w(0) or do_read_nonvolatile;
	wire_w_lg_w_lg_w_lg_do_sec_erase532w533w534w(0) <= wire_w_lg_w_lg_do_sec_erase532w533w(0) or do_die_erase;
	wire_w_lg_w_lg_w_lg_do_write72w116w117w(0) <= wire_w_lg_w_lg_do_write72w116w(0) or do_die_erase;
	wire_w_lg_w_lg_bp3_wire539w540w(0) <= wire_w_lg_bp3_wire539w(0) or bp1_wire;
	wire_w_lg_w_lg_do_read407w442w(0) <= wire_w_lg_do_read407w(0) or do_read_sid;
	wire_w_lg_w_lg_do_read407w428w(0) <= wire_w_lg_do_read407w(0) or do_write;
	wire_w_lg_w_lg_do_read_sid147w148w(0) <= wire_w_lg_do_read_sid147w(0) or do_sec_erase;
	wire_w_lg_w_lg_do_read_stat438w439w(0) <= wire_w_lg_do_read_stat438w(0) or do_read_volatile;
	wire_w_lg_w_lg_do_sec_erase532w533w(0) <= wire_w_lg_do_sec_erase532w(0) or do_bulk_erase;
	wire_w_lg_w_lg_do_write72w116w(0) <= wire_w_lg_do_write72w(0) or do_bulk_erase;
	wire_w_lg_w_lg_do_write72w73w(0) <= wire_w_lg_do_write72w(0) or do_die_erase;
	wire_w_lg_w_lg_w_prot_wire_range551w570w572w(0) <= wire_w_lg_w_prot_wire_range551w570w(0) or wire_w_prot_wire_range556w(0);
	wire_w_lg_bp3_wire539w(0) <= bp3_wire or bp2_wire;
	wire_w_lg_data0out_wire446w(0) <= data0out_wire or wire_w_dataout_wire_range445w(0);
	wire_w_lg_do_4baddr341w(0) <= do_4baddr or wire_w_lg_do_ex4baddr340w(0);
	wire_w_lg_do_ex4baddr340w(0) <= do_ex4baddr or wire_w_lg_do_bulk_erase339w(0);
	wire_w_lg_do_read407w(0) <= do_read or do_fast_read;
	wire_w_lg_do_read_rdid125w(0) <= do_read_rdid or wire_w_lg_w_lg_do_read_stat123w124w(0);
	wire_w_lg_do_read_sid147w(0) <= do_read_sid or do_write;
	wire_w_lg_do_read_stat438w(0) <= do_read_stat or do_read_rdid;
	wire_w_lg_do_sec_erase54w(0) <= do_sec_erase or do_die_erase;
	wire_w_lg_do_sec_erase532w(0) <= do_sec_erase or do_write;
	wire_w_lg_do_wren342w(0) <= do_wren or wire_w_lg_do_4baddr341w(0);
	wire_w_lg_do_write72w(0) <= do_write or do_sec_erase;
	wire_w_lg_end_operation502w(0) <= end_operation or wire_w_lg_w_lg_do_polling500w501w(0);
	wire_w_lg_load_opcode315w(0) <= load_opcode or shift_opcode;
	wire_w_lg_rden_wire412w(0) <= rden_wire or wren_wire;
	wire_w_lg_w_mask_prot_add_range583w597w(0) <= wire_w_mask_prot_add_range583w(0) or wire_w_mask_prot_comp_tb_range593w(0);
	wire_w_lg_w_mask_prot_add_range588w601w(0) <= wire_w_mask_prot_add_range588w(0) or wire_w_mask_prot_comp_tb_range598w(0);
	wire_w_lg_w_mask_prot_check_range585w595w(0) <= wire_w_mask_prot_check_range585w(0) or wire_w_mask_prot_comp_ntb_range591w(0);
	wire_w_lg_w_mask_prot_check_range590w599w(0) <= wire_w_mask_prot_check_range590w(0) or wire_w_mask_prot_comp_ntb_range596w(0);
	wire_w_lg_w_prot_wire_range551w570w(0) <= wire_w_prot_wire_range551w(0) or wire_w_prot_wire_range553w(0);
	wire_w_lg_w_mask_prot_range568w578w(0) <= wire_w_mask_prot_range568w(0) xor wire_w_mask_prot_add_range576w(0);
	wire_w_lg_w_mask_prot_range571w584w(0) <= wire_w_mask_prot_range571w(0) xor wire_w_mask_prot_add_range583w(0);
	wire_w_lg_w_mask_prot_range573w589w(0) <= wire_w_mask_prot_range573w(0) xor wire_w_mask_prot_add_range588w(0);
	addr_overdie <= '0';
	addr_overdie_pos <= '0';
	addr_reg_overdie <= (others => '0');
	b4addr_opcode <= (others => '0');
	be_write_prot <= ((do_bulk_erase or do_die_erase) and wire_w_lg_w_lg_w_lg_bp3_wire539w540w541w(0));
	berase_opcode <= (others => '0');
	bp0_wire <= statreg_int(2);
	bp1_wire <= statreg_int(3);
	bp2_wire <= statreg_int(4);
	bp3_wire <= statreg_int(6);
	busy <= busy_wire;
	busy_wire <= ((((((((((((((do_read_rdid or do_read_sid) or do_read) or do_fast_read) or do_write) or do_sec_prot) or do_read_stat) or do_sec_erase) or do_bulk_erase) or do_die_erase) or do_4baddr) or do_read_volatile) or do_fread_epcq) or do_read_nonvolatile) or do_ex4baddr);
	clkin_wire <= clkin;
	clr_addmsb_wire <= ((wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range103w108w420w421w(0) or wire_w_lg_w_lg_w_lg_do_read359w360w419w(0)) or wire_w_lg_w_lg_w_lg_w_lg_do_sec_erase54w416w417w418w(0));
	clr_endrbyte_wire <= ((((wire_w_lg_do_read407w(0) and (not wire_gen_cntr_q(2))) and wire_gen_cntr_q(1)) and wire_gen_cntr_q(0)) or clr_read_wire2);
	clr_read_wire <= clr_read_reg;
	clr_read_wire2 <= clr_read_reg2;
	clr_rstat_wire <= clr_rstat_reg;
	clr_write_wire <= clr_write_reg;
	clr_write_wire2 <= clr_write_reg2;
	data0out_wire <= wire_cycloneii_asmiblock2_data0out;
	data_valid <= data_valid_wire;
	data_valid_wire <= dvalid_reg2;
	datain_reg_wire_in <= ( wire_w_lg_w_lg_not_busy617w618w & wire_w_lg_not_busy622w);
	datain_wire <= ( "0000");
	dataout <= ( read_data_reg(7 downto 0));
	dataout_wire <= ( "0000");
	derase_opcode <= (others => '0');
	do_4baddr <= '0';
	do_bulk_erase <= '0';
	do_die_erase <= '0';
	do_ex4baddr <= '0';
	do_fast_read <= '0';
	do_fread_epcq <= '0';
	do_freadwrv_polling <= '0';
	do_memadd <= do_wrmemadd_reg;
	do_polling <= ((do_write_polling or do_sprot_polling) or do_freadwrv_polling);
	do_read <= (((wire_w_lg_read_rdid_wire9w(0) and wire_w_lg_read_sid_wire8w(0)) and wire_w_lg_sec_protect_wire7w(0)) and read_wire);
	do_read_nonvolatile <= '0';
	do_read_rdid <= '0';
	do_read_sid <= '0';
	do_read_stat <= ((((((((wire_w_lg_read_rdid_wire9w(0) and wire_w_lg_read_sid_wire8w(0)) and wire_w_lg_sec_protect_wire7w(0)) and (not (read_wire or fast_read_wire))) and wire_w_lg_write_wire17w(0)) and read_status_wire) or do_write_rstat) or do_sprot_rstat) or do_write_volatile_rstat);
	do_read_volatile <= '0';
	do_sec_erase <= '0';
	do_sec_prot <= '0';
	do_secprot_wren <= '0';
	do_sprot_polling <= '0';
	do_sprot_rstat <= '0';
	do_wait_dummyclk <= '0';
	do_wren <= ((do_write_wren or do_secprot_wren) or do_write_volatile_wren);
	do_write <= ((((wire_w_lg_read_rdid_wire9w(0) and wire_w_lg_read_sid_wire8w(0)) and wire_w_lg_sec_protect_wire7w(0)) and (not (read_wire or fast_read_wire))) and write_wire);
	do_write_polling <= wire_w_lg_w_lg_w530w641w642w(0);
	do_write_rstat <= write_rstat_reg;
	do_write_volatile <= '0';
	do_write_volatile_rstat <= '0';
	do_write_volatile_wren <= '0';
	do_write_wren <= ((not wire_wrstage_cntr_q(1)) and wire_wrstage_cntr_q(0));
	end1_cyc_gen_cntr_wire <= (wire_gen_cntr_w_lg_w_q_range113w114w(0) and (not wire_gen_cntr_q(0)));
	end1_cyc_normal_in_wire <= ((((((((((wire_stage_cntr_w_lg_w_lg_w_q_range102w107w133w(0) and (not wire_gen_cntr_q(2))) and wire_gen_cntr_q(1)) and wire_gen_cntr_q(0)) or wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range102w107w133w134w135w(0)) or (do_read and end_read)) or (do_fast_read and end_fast_read)) or wire_w_lg_w_lg_w_lg_w_lg_do_write72w116w117w130w(0)) or wire_w_lg_do_write70w(0)) or ((do_read_stat and start_poll) and wire_w_lg_st_busy_wire127w(0))) or wire_w_lg_w_lg_do_read_rdid125w126w(0));
	end1_cyc_reg_in_wire <= end1_cyc_normal_in_wire;
	end_add_cycle <= wire_mux211_dataout;
	end_add_cycle_mux_datab_wire <= (wire_addbyte_cntr_q(2) and wire_addbyte_cntr_q(1));
	end_fast_read <= end_read_reg;
	end_one_cyc_pos <= end1_cyc_reg2;
	end_one_cycle <= end1_cyc_reg;
	end_op_wire <= (((((((((((wire_stage_cntr_w_lg_w_q_range103w108w(0) and ((wire_w_lg_w_lg_w_lg_w_lg_do_read359w360w361w362w(0) or (do_read and end_read)) or (do_fast_read and end_fast_read))) or (wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range103w106w354w355w(0) and wire_w_lg_do_polling203w(0))) or ((((((do_read_rdid and end_one_cyc_pos) and wire_stage_cntr_q(1)) and wire_stage_cntr_q(0)) and wire_addbyte_cntr_q(2)) and wire_addbyte_cntr_q(1)) and wire_addbyte_cntr_w_lg_w_q_range161w162w(0))) or (wire_w_lg_w_lg_start_poll345w346w(0) and wire_w_lg_st_busy_wire127w(0))) or wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range103w104w105w343w344w(0)) or wire_w_lg_w_lg_w_lg_w_lg_do_write72w116w117w130w(0)) or wire_w_lg_w_lg_do_write63w338w(0)) or wire_w_lg_do_write70w(0)) or wire_stage_cntr_w337w(0)) or wire_stage_cntr_w_lg_w332w333w(0)) or (wire_stage_cntr_w_lg_w_lg_w_q_range103w106w327w(0) and ((do_write_volatile or do_read_volatile) or wire_w_lg_do_read_nonvolatile325w(0))));
	end_operation <= end_op_reg;
	end_ophdly <= end_op_hdlyreg;
	end_pgwr_data <= '0';
	end_read <= end_read_reg;
	end_read_byte <= (end_rbyte_reg and wire_w_lg_addr_overdie490w(0));
	end_wrstage <= end_operation;
	exb4addr_opcode <= (others => '0');
	fast_read_opcode <= (others => '0');
	fast_read_wire <= '0';
	freadwrv_sdoin <= '0';
	ill_write_wire <= ill_write_reg;
	illegal_write <= ill_write_wire;
	illegal_write_b4out_wire <= (((do_write and write_prot_true) or (illegal_write_prot and write_prot_true2)) or wire_w_lg_do_write70w(0));
	illegal_write_prot <= illegal_write_prot_reg;
	in_operation <= busy_wire;
	load_opcode <= ((((wire_stage_cntr_w_lg_w_q_range103w104w(0) and wire_stage_cntr_w_lg_w_q_range102w107w(0)) and (not wire_gen_cntr_q(2))) and wire_gen_cntr_w_lg_w_q_range111w112w(0)) and wire_gen_cntr_q(0));
	mask_prot <= ( wire_w_lg_w_lg_w_prot_wire_range551w570w572w & wire_w_lg_w_prot_wire_range551w570w & prot_wire(1));
	mask_prot_add <= ( wire_w_lg_w_mask_prot_range573w587w & wire_w_lg_w_mask_prot_range571w582w & wire_w_lg_w_mask_prot_range568w575w);
	mask_prot_check <= ( wire_w_lg_w_mask_prot_range573w589w & wire_w_lg_w_mask_prot_range571w584w & wire_w_lg_w_mask_prot_range568w578w);
	mask_prot_comp_ntb <= ( wire_w_lg_w_mask_prot_check_range590w599w & wire_w_lg_w_mask_prot_check_range585w595w & mask_prot_check(0));
	mask_prot_comp_tb <= ( wire_w_lg_w_mask_prot_add_range588w601w & wire_w_lg_w_mask_prot_add_range583w597w & mask_prot_add(0));
	memadd_sdoin <= add_msb_reg;
	ncs_reg_ena_wire <= (((wire_stage_cntr_w_lg_w_lg_w_q_range103w104w105w(0) and end_one_cyc_pos) or addr_overdie_pos) or end_operation);
	not_busy <= busy_det_reg;
	oe_wire <= '0';
	pagewr_buf_not_empty <= ( "1");
	prot_wire <= ( wire_w_lg_w_lg_bp2_wire564w567w & wire_w_lg_w_lg_bp2_wire564w565w & wire_w_lg_w_lg_bp2_wire559w562w & wire_w_lg_w_lg_bp2_wire559w560w & wire_w_lg_w_lg_w_lg_bp2_wire547w554w557w & wire_w_lg_w_lg_w_lg_bp2_wire547w554w555w & wire_w_lg_w_lg_w_lg_bp2_wire547w548w552w & wire_w_lg_w_lg_w_lg_bp2_wire547w548w549w);
	rden_wire <= rden;
	rdid_opcode <= (others => '0');
	rdummyclk_opcode <= (others => '0');
	read_data_reg_in_wire <= ( read_dout_reg(7 downto 0));
	read_opcode <= "00000011";
	read_rdid_wire <= '0';
	read_sid_wire <= '0';
	read_status_wire <= '0';
	read_wire <= read_reg;
	rflagstat_opcode <= "00000101";
	rnvdummyclk_opcode <= (others => '0');
	rsid_opcode <= (others => '0');
	rsid_sdoin <= '0';
	rstat_opcode <= "00000101";
	scein_wire <= wire_ncs_reg_w_lg_q380w(0);
	sdoin_wire <= to_sdoin_wire;
	sec_protect_wire <= '0';
	secprot_opcode <= (others => '0');
	secprot_sdoin <= '0';
	serase_opcode <= (others => '0');
	shift_opcode <= shift_op_reg;
	shift_opdata <= stage2_wire;
	shift_pgwr_data <= '0';
	st_busy_wire <= statreg_int(0);
	stage2_wire <= stage2_reg;
	stage3_wire <= stage3_reg;
	stage4_wire <= stage4_reg;
	start_frpoll <= '0';
	start_poll <= ((start_wrpoll or start_sppoll) or start_frpoll);
	start_sppoll <= '0';
	start_wrpoll <= start_wrpoll_reg2;
	to_sdoin_wire <= ((((((shift_opdata and asmi_opcode_reg(7)) or rsid_sdoin) or memadd_sdoin) or write_sdoin) or secprot_sdoin) or freadwrv_sdoin);
	wren_opcode <= "00000110";
	wren_wire <= wren;
	write_opcode <= "00000010";
	write_prot_true <= write_prot_reg;
	write_prot_true2 <= write_prot_reg2;
	write_sdoin <= ((((do_write and stage4_wire) and wire_wrstage_cntr_q(1)) and wire_wrstage_cntr_q(0)) and wrsdoin_reg);
	write_wire <= write_reg;
	wrvolatile_opcode <= (others => '0');
	wire_w_addr_range403w(0) <= addr(0);
	wire_w_addr_range395w <= addr(23 downto 1);
	wire_w_addr_reg_overdie_range401w(0) <= addr_reg_overdie(0);
	wire_w_addr_reg_overdie_range391w <= addr_reg_overdie(23 downto 1);
	wire_w_b4addr_opcode_range266w(0) <= b4addr_opcode(0);
	wire_w_b4addr_opcode_range175w <= b4addr_opcode(7 downto 1);
	wire_w_berase_opcode_range270w(0) <= berase_opcode(0);
	wire_w_berase_opcode_range183w <= berase_opcode(7 downto 1);
	wire_w_datain_range621w(0) <= datain(0);
	wire_w_datain_range616w <= datain(7 downto 1);
	wire_w_dataout_wire_range445w(0) <= dataout_wire(1);
	wire_w_derase_opcode_range272w(0) <= derase_opcode(0);
	wire_w_derase_opcode_range188w <= derase_opcode(7 downto 1);
	wire_w_exb4addr_opcode_range264w(0) <= exb4addr_opcode(0);
	wire_w_exb4addr_opcode_range170w <= exb4addr_opcode(7 downto 1);
	wire_w_fast_read_opcode_range288w(0) <= fast_read_opcode(0);
	wire_w_fast_read_opcode_range228w <= fast_read_opcode(7 downto 1);
	wire_w_mask_prot_range568w(0) <= mask_prot(0);
	wire_w_mask_prot_range571w(0) <= mask_prot(1);
	wire_w_mask_prot_range573w(0) <= mask_prot(2);
	wire_w_mask_prot_add_range576w(0) <= mask_prot_add(0);
	wire_w_mask_prot_add_range583w(0) <= mask_prot_add(1);
	wire_w_mask_prot_add_range588w(0) <= mask_prot_add(2);
	wire_w_mask_prot_check_range585w(0) <= mask_prot_check(1);
	wire_w_mask_prot_check_range590w(0) <= mask_prot_check(2);
	wire_w_mask_prot_comp_ntb_range591w(0) <= mask_prot_comp_ntb(0);
	wire_w_mask_prot_comp_ntb_range596w(0) <= mask_prot_comp_ntb(1);
	wire_w_mask_prot_comp_tb_range593w(0) <= mask_prot_comp_tb(0);
	wire_w_mask_prot_comp_tb_range598w(0) <= mask_prot_comp_tb(1);
	wire_w_pagewr_buf_not_empty_range68w(0) <= pagewr_buf_not_empty(0);
	wire_w_prot_wire_range551w(0) <= prot_wire(1);
	wire_w_prot_wire_range553w(0) <= prot_wire(2);
	wire_w_prot_wire_range556w(0) <= prot_wire(3);
	wire_w_rdid_opcode_range294w(0) <= rdid_opcode(0);
	wire_w_rdid_opcode_range239w <= rdid_opcode(7 downto 1);
	wire_w_rdummyclk_opcode_range286w(0) <= rdummyclk_opcode(0);
	wire_w_rdummyclk_opcode_range221w <= rdummyclk_opcode(7 downto 1);
	wire_w_read_opcode_range290w(0) <= read_opcode(0);
	wire_w_read_opcode_range231w <= read_opcode(7 downto 1);
	wire_w_rflagstat_opcode_range276w(0) <= rflagstat_opcode(0);
	wire_w_rflagstat_opcode_range198w <= rflagstat_opcode(7 downto 1);
	wire_w_rnvdummyclk_opcode_range282w(0) <= rnvdummyclk_opcode(0);
	wire_w_rnvdummyclk_opcode_range211w <= rnvdummyclk_opcode(7 downto 1);
	wire_w_rsid_opcode_range296w(0) <= rsid_opcode(0);
	wire_w_rsid_opcode_range242w <= rsid_opcode(7 downto 1);
	wire_w_rstat_opcode_range278w(0) <= rstat_opcode(0);
	wire_w_rstat_opcode_range202w <= rstat_opcode(7 downto 1);
	wire_w_secprot_opcode_range292w(0) <= secprot_opcode(0);
	wire_w_secprot_opcode_range234w <= secprot_opcode(7 downto 1);
	wire_w_serase_opcode_range274w(0) <= serase_opcode(0);
	wire_w_serase_opcode_range193w <= serase_opcode(7 downto 1);
	wire_w_wren_opcode_range268w(0) <= wren_opcode(0);
	wire_w_wren_opcode_range180w <= wren_opcode(7 downto 1);
	wire_w_write_opcode_range280w(0) <= write_opcode(0);
	wire_w_write_opcode_range206w <= write_opcode(7 downto 1);
	wire_w_wrvolatile_opcode_range284w(0) <= wrvolatile_opcode(0);
	wire_w_wrvolatile_opcode_range214w <= wrvolatile_opcode(7 downto 1);
	wire_addbyte_cntr_w_lg_w_q_range158w163w(0) <= wire_addbyte_cntr_w_q_range158w(0) and wire_addbyte_cntr_w_lg_w_q_range161w162w(0);
	wire_addbyte_cntr_w_lg_w_q_range161w162w(0) <= not wire_addbyte_cntr_w_q_range161w(0);
	wire_addbyte_cntr_clk_en <= wire_stage_cntr_w157w(0);
	wire_stage_cntr_w157w(0) <= ((wire_stage_cntr_w_lg_w_lg_w_q_range103w106w154w(0) and wire_w_lg_w_lg_w151w152w153w(0)) or addr_overdie) or end_operation;
	wire_addbyte_cntr_clock <= wire_w_lg_clkin_wire101w(0);
	wire_addbyte_cntr_sclr <= wire_w_lg_end_operation100w(0);
	wire_w_lg_end_operation100w(0) <= end_operation or addr_overdie;
	wire_addbyte_cntr_w_q_range161w(0) <= wire_addbyte_cntr_q(0);
	wire_addbyte_cntr_w_q_range158w(0) <= wire_addbyte_cntr_q(1);
	addbyte_cntr :  a_graycounter
	  generic map (
		width => 3
	  )
	  port map ( 
		aclr => reset,
		clk_en => wire_addbyte_cntr_clk_en,
		clock => wire_addbyte_cntr_clock,
		q => wire_addbyte_cntr_q,
		sclr => wire_addbyte_cntr_sclr
	  );
	wire_gen_cntr_w_lg_w_q_range113w114w(0) <= wire_gen_cntr_w_q_range113w(0) and wire_gen_cntr_w_lg_w_q_range111w112w(0);
	wire_gen_cntr_w_lg_w_q_range111w112w(0) <= not wire_gen_cntr_w_q_range111w(0);
	wire_gen_cntr_clk_en <= wire_w_lg_w_lg_w_lg_in_operation40w41w42w(0);
	wire_w_lg_w_lg_w_lg_in_operation40w41w42w(0) <= ((in_operation and wire_w_lg_end_ophdly39w(0)) or do_wait_dummyclk) or addr_overdie;
	wire_gen_cntr_sclr <= wire_w_lg_w_lg_end1_cyc_reg_in_wire43w44w(0);
	wire_w_lg_w_lg_end1_cyc_reg_in_wire43w44w(0) <= (end1_cyc_reg_in_wire or addr_overdie) or do_wait_dummyclk;
	wire_gen_cntr_w_q_range111w(0) <= wire_gen_cntr_q(1);
	wire_gen_cntr_w_q_range113w(0) <= wire_gen_cntr_q(2);
	gen_cntr :  a_graycounter
	  generic map (
		width => 3
	  )
	  port map ( 
		aclr => reset,
		clk_en => wire_gen_cntr_clk_en,
		clock => clkin_wire,
		q => wire_gen_cntr_q,
		sclr => wire_gen_cntr_sclr
	  );
	wire_stage_cntr_w_lg_w332w333w(0) <= wire_stage_cntr_w332w(0) and end_one_cycle;
	wire_stage_cntr_w332w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range103w106w329w330w331w(0) and end_add_cycle;
	wire_stage_cntr_w337w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range103w106w334w335w336w(0) and end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range103w106w329w330w331w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range103w106w329w330w(0) and wire_w_lg_do_read_stat52w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range103w106w334w335w336w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range103w106w334w335w(0) and wire_w_lg_do_read_stat52w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range103w104w105w343w344w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range103w104w105w343w(0) and end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range103w108w420w421w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range103w108w420w(0) and end_one_cyc_pos;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range103w106w329w330w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range103w106w329w(0) and wire_w_lg_do_wren53w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range103w106w354w355w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range103w106w354w(0) and end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range103w106w334w335w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range103w106w334w(0) and wire_w_lg_do_wren53w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range103w104w105w343w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range103w104w105w(0) and wire_w_lg_do_wren342w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range103w108w420w(0) <= wire_stage_cntr_w_lg_w_q_range103w108w(0) and end_add_cycle;
	wire_stage_cntr_w_lg_w_lg_w_q_range103w106w329w(0) <= wire_stage_cntr_w_lg_w_q_range103w106w(0) and wire_w_lg_do_sec_erase54w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range103w106w354w(0) <= wire_stage_cntr_w_lg_w_q_range103w106w(0) and do_read_stat;
	wire_stage_cntr_w_lg_w_lg_w_q_range103w106w334w(0) <= wire_stage_cntr_w_lg_w_q_range103w106w(0) and do_sec_prot;
	wire_stage_cntr_w_lg_w_lg_w_q_range103w106w154w(0) <= wire_stage_cntr_w_lg_w_q_range103w106w(0) and end_one_cyc_pos;
	wire_stage_cntr_w_lg_w_lg_w_q_range103w106w327w(0) <= wire_stage_cntr_w_lg_w_q_range103w106w(0) and end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range102w107w133w134w135w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range102w107w133w134w(0) and end1_cyc_gen_cntr_wire;
	wire_stage_cntr_w_lg_w_lg_w_q_range102w107w133w(0) <= wire_stage_cntr_w_lg_w_q_range102w107w(0) and wire_stage_cntr_w_lg_w_q_range103w104w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range103w104w105w(0) <= wire_stage_cntr_w_lg_w_q_range103w104w(0) and wire_stage_cntr_w_q_range102w(0);
	wire_stage_cntr_w_lg_w_q_range103w108w(0) <= wire_stage_cntr_w_q_range103w(0) and wire_stage_cntr_w_lg_w_q_range102w107w(0);
	wire_stage_cntr_w_lg_w_q_range103w106w(0) <= wire_stage_cntr_w_q_range103w(0) and wire_stage_cntr_w_q_range102w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range102w107w133w134w(0) <= not wire_stage_cntr_w_lg_w_lg_w_q_range102w107w133w(0);
	wire_stage_cntr_w_lg_w_q_range102w107w(0) <= not wire_stage_cntr_w_q_range102w(0);
	wire_stage_cntr_w_lg_w_q_range103w104w(0) <= not wire_stage_cntr_w_q_range103w(0);
	wire_stage_cntr_clk_en <= wire_w_lg_w_lg_w_lg_w96w97w98w99w(0);
	wire_w_lg_w_lg_w_lg_w96w97w98w99w(0) <= (((((((((((((in_operation and end_one_cycle) and (not (stage3_wire and wire_w_lg_end_add_cycle83w(0)))) and (not (stage4_wire and wire_w_lg_end_read80w(0)))) and (not (stage4_wire and wire_w_lg_end_fast_read77w(0)))) and (not ((wire_w_lg_w_lg_do_write72w73w(0) or do_bulk_erase) and write_prot_true))) and (not wire_w_lg_do_write70w(0))) and (not (stage3_wire and st_busy_wire))) and (not (wire_w_lg_do_write63w(0) and wire_w_lg_end_pgwr_data62w(0)))) and (not (stage2_wire and do_wren))) and (not (((wire_w_lg_stage3_wire55w(0) and wire_w_lg_do_wren53w(0)) and wire_w_lg_do_read_stat52w(0)) and wire_w_lg_do_read_rdid51w(0)))) and (not (stage3_wire and ((do_write_volatile or do_read_volatile) or do_read_nonvolatile)))) or wire_w_lg_w_lg_stage3_wire45w46w(0)) or addr_overdie) or end_ophdly;
	wire_stage_cntr_sclr <= wire_w_lg_end_operation100w(0);
	wire_stage_cntr_w_q_range102w(0) <= wire_stage_cntr_q(0);
	wire_stage_cntr_w_q_range103w(0) <= wire_stage_cntr_q(1);
	stage_cntr :  a_graycounter
	  generic map (
		width => 2
	  )
	  port map ( 
		aclr => reset,
		clk_en => wire_stage_cntr_clk_en,
		clock => clkin_wire,
		q => wire_stage_cntr_q,
		sclr => wire_stage_cntr_sclr
	  );
	wire_wrstage_cntr_w_lg_w_q_range524w525w(0) <= wire_wrstage_cntr_w_q_range524w(0) and wire_wrstage_cntr_w_lg_w_q_range522w523w(0);
	wire_wrstage_cntr_w_lg_w_q_range522w523w(0) <= not wire_wrstage_cntr_w_q_range522w(0);
	wire_wrstage_cntr_clk_en <= wire_w_lg_w_lg_w_lg_w_lg_w517w518w519w520w521w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w517w518w519w520w521w(0) <= (wire_w_lg_w_lg_w517w518w519w(0) and wire_w_lg_st_busy_wire127w(0)) or clr_write_wire2;
	wire_wrstage_cntr_clock <= wire_w_lg_clkin_wire101w(0);
	wire_wrstage_cntr_w_q_range522w(0) <= wire_wrstage_cntr_q(0);
	wire_wrstage_cntr_w_q_range524w(0) <= wire_wrstage_cntr_q(1);
	wrstage_cntr :  a_graycounter
	  generic map (
		width => 2
	  )
	  port map ( 
		aclr => reset,
		clk_en => wire_wrstage_cntr_clk_en,
		clock => wire_wrstage_cntr_clock,
		q => wire_wrstage_cntr_q,
		sclr => clr_write_wire2
	  );
	wire_cycloneii_asmiblock2_sdoin <= wire_w_lg_sdoin_wire320w(0);
	wire_w_lg_sdoin_wire320w(0) <= sdoin_wire or datain_wire(0);
	cycloneii_asmiblock2 :  cycloneii_asmiblock
	  port map ( 
		data0out => wire_cycloneii_asmiblock2_data0out,
		dclkin => clkin_wire,
		oe => oe_wire,
		scein => scein_wire,
		sdoin => wire_cycloneii_asmiblock2_sdoin
	  );
	process (clkin_wire, reset)
	begin
		if (reset = '1') then add_msb_reg <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then 
			if (wire_add_msb_reg_ena = '1') then 
				if (clr_addmsb_wire = '1') then add_msb_reg <= '0';
				else add_msb_reg <= addr_reg(23);
				end if;
			end if;
		end if;
	end process;
	wire_add_msb_reg_ena <= ((((wire_w_lg_w_lg_w_lg_w_lg_do_read407w428w429w430w(0) and (not (wire_w_lg_w_lg_do_write72w73w(0) and wire_w_lg_do_memadd425w(0)))) and wire_stage_cntr_q(1)) and wire_stage_cntr_q(0)) or clr_addmsb_wire);
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(0) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(0) = '1') then addr_reg(0) <= wire_addr_reg_d(0);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(1) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(1) = '1') then addr_reg(1) <= wire_addr_reg_d(1);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(2) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(2) = '1') then addr_reg(2) <= wire_addr_reg_d(2);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(3) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(3) = '1') then addr_reg(3) <= wire_addr_reg_d(3);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(4) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(4) = '1') then addr_reg(4) <= wire_addr_reg_d(4);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(5) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(5) = '1') then addr_reg(5) <= wire_addr_reg_d(5);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(6) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(6) = '1') then addr_reg(6) <= wire_addr_reg_d(6);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(7) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(7) = '1') then addr_reg(7) <= wire_addr_reg_d(7);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(8) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(8) = '1') then addr_reg(8) <= wire_addr_reg_d(8);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(9) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(9) = '1') then addr_reg(9) <= wire_addr_reg_d(9);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(10) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(10) = '1') then addr_reg(10) <= wire_addr_reg_d(10);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(11) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(11) = '1') then addr_reg(11) <= wire_addr_reg_d(11);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(12) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(12) = '1') then addr_reg(12) <= wire_addr_reg_d(12);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(13) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(13) = '1') then addr_reg(13) <= wire_addr_reg_d(13);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(14) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(14) = '1') then addr_reg(14) <= wire_addr_reg_d(14);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(15) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(15) = '1') then addr_reg(15) <= wire_addr_reg_d(15);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(16) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(16) = '1') then addr_reg(16) <= wire_addr_reg_d(16);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(17) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(17) = '1') then addr_reg(17) <= wire_addr_reg_d(17);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(18) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(18) = '1') then addr_reg(18) <= wire_addr_reg_d(18);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(19) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(19) = '1') then addr_reg(19) <= wire_addr_reg_d(19);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(20) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(20) = '1') then addr_reg(20) <= wire_addr_reg_d(20);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(21) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(21) = '1') then addr_reg(21) <= wire_addr_reg_d(21);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(22) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(22) = '1') then addr_reg(22) <= wire_addr_reg_d(22);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then addr_reg(23) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_addr_reg_ena(23) = '1') then addr_reg(23) <= wire_addr_reg_d(23);
			end if;
		end if;
	end process;
	wire_addr_reg_d <= ( wire_w_lg_w_lg_w_lg_not_busy396w397w398w & wire_w_lg_w_lg_not_busy404w405w);
	loop43 : for i in 0 to 23 generate
		wire_addr_reg_ena(i) <= wire_w_lg_w_lg_w_lg_w_lg_rden_wire412w413w414w415w(0);
	end generate loop43;
	wire_addr_reg_w_q_range574w(0) <= addr_reg(16);
	wire_addr_reg_w_q_range581w(0) <= addr_reg(17);
	wire_addr_reg_w_q_range393w <= addr_reg(22 downto 0);
	wire_addr_reg_w_q_range586w(0) <= addr_reg(18);
	process (clkin_wire, reset)
	begin
		if (reset = '1') then asmi_opcode_reg(0) <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then 
			if (wire_asmi_opcode_reg_ena(0) = '1') then asmi_opcode_reg(0) <= wire_asmi_opcode_reg_d(0);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then asmi_opcode_reg(1) <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then 
			if (wire_asmi_opcode_reg_ena(1) = '1') then asmi_opcode_reg(1) <= wire_asmi_opcode_reg_d(1);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then asmi_opcode_reg(2) <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then 
			if (wire_asmi_opcode_reg_ena(2) = '1') then asmi_opcode_reg(2) <= wire_asmi_opcode_reg_d(2);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then asmi_opcode_reg(3) <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then 
			if (wire_asmi_opcode_reg_ena(3) = '1') then asmi_opcode_reg(3) <= wire_asmi_opcode_reg_d(3);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then asmi_opcode_reg(4) <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then 
			if (wire_asmi_opcode_reg_ena(4) = '1') then asmi_opcode_reg(4) <= wire_asmi_opcode_reg_d(4);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then asmi_opcode_reg(5) <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then 
			if (wire_asmi_opcode_reg_ena(5) = '1') then asmi_opcode_reg(5) <= wire_asmi_opcode_reg_d(5);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then asmi_opcode_reg(6) <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then 
			if (wire_asmi_opcode_reg_ena(6) = '1') then asmi_opcode_reg(6) <= wire_asmi_opcode_reg_d(6);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then asmi_opcode_reg(7) <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then 
			if (wire_asmi_opcode_reg_ena(7) = '1') then asmi_opcode_reg(7) <= wire_asmi_opcode_reg_d(7);
			end if;
		end if;
	end process;
	wire_asmi_opcode_reg_d <= ( wire_w_lg_w_lg_w259w260w261w & wire_w_lg_w312w313w);
	loop44 : for i in 0 to 7 generate
		wire_asmi_opcode_reg_ena(i) <= wire_w_lg_load_opcode315w(0);
	end generate loop44;
	wire_asmi_opcode_reg_w_q_range168w <= asmi_opcode_reg(6 downto 0);
	process (clkin_wire, reset)
	begin
		if (reset = '1') then busy_det_reg <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then busy_det_reg <= wire_w_lg_busy_wire1w(0);
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then clr_read_reg <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then clr_read_reg <= ((do_read_sid or do_sec_prot) or end_operation);
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then clr_read_reg2 <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then clr_read_reg2 <= clr_read_reg;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then clr_rstat_reg <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then clr_rstat_reg <= ((end_operation or do_read_sid) or do_read);
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then clr_write_reg <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then clr_write_reg <= ((((((wire_w_lg_w_lg_w_lg_w_lg_w530w641w642w658w659w(0) or wire_w_lg_do_write70w(0)) or wire_w_lg_w_lg_w655w656w657w(0)) or do_read_sid) or do_sec_prot) or do_read) or do_fast_read);
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then clr_write_reg2 <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then clr_write_reg2 <= clr_write_reg;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then datain_reg(0) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_datain_reg_ena(0) = '1') then datain_reg(0) <= wire_datain_reg_d(0);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then datain_reg(1) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_datain_reg_ena(1) = '1') then datain_reg(1) <= wire_datain_reg_d(1);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then datain_reg(2) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_datain_reg_ena(2) = '1') then datain_reg(2) <= wire_datain_reg_d(2);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then datain_reg(3) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_datain_reg_ena(3) = '1') then datain_reg(3) <= wire_datain_reg_d(3);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then datain_reg(4) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_datain_reg_ena(4) = '1') then datain_reg(4) <= wire_datain_reg_d(4);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then datain_reg(5) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_datain_reg_ena(5) = '1') then datain_reg(5) <= wire_datain_reg_d(5);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then datain_reg(6) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_datain_reg_ena(6) = '1') then datain_reg(6) <= wire_datain_reg_d(6);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then datain_reg(7) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_datain_reg_ena(7) = '1') then datain_reg(7) <= wire_datain_reg_d(7);
			end if;
		end if;
	end process;
	wire_datain_reg_d <= ( datain_reg_wire_in(7 downto 0));
	loop45 : for i in 0 to 7 generate
		wire_datain_reg_ena(i) <= wire_w_lg_w_lg_wren_wire631w632w(0);
	end generate loop45;
	wire_datain_reg_w_q_range614w <= datain_reg(6 downto 0);
	process (clkin_wire, reset)
	begin
		if (reset = '1') then do_wrmemadd_reg <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then do_wrmemadd_reg <= (wire_wrstage_cntr_q(1) and wire_wrstage_cntr_q(0));
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then dvalid_reg <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_dvalid_reg_ena = '1') then 
				if (wire_dvalid_reg_sclr = '1') then dvalid_reg <= '0';
				else dvalid_reg <= (end_read_byte and end_one_cyc_pos);
				end if;
			end if;
		end if;
	end process;
	wire_dvalid_reg_ena <= wire_w_lg_do_read407w(0);
	wire_dvalid_reg_sclr <= (end_op_wire or end_operation);
	process (clkin_wire, reset)
	begin
		if (reset = '1') then dvalid_reg2 <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then dvalid_reg2 <= dvalid_reg;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then end1_cyc_reg <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then end1_cyc_reg <= end1_cyc_reg_in_wire;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then end1_cyc_reg2 <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then end1_cyc_reg2 <= end_one_cycle;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then end_op_hdlyreg <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then end_op_hdlyreg <= end_operation;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then end_op_reg <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then end_op_reg <= end_op_wire;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then end_rbyte_reg <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_end_rbyte_reg_ena = '1') then 
				if (wire_end_rbyte_reg_sclr = '1') then end_rbyte_reg <= '0';
				else end_rbyte_reg <= wire_w_lg_w_lg_w_lg_do_read407w474w475w(0);
				end if;
			end if;
		end if;
	end process;
	wire_end_rbyte_reg_ena <= ((wire_gen_cntr_w_lg_w_q_range113w114w(0) and wire_gen_cntr_q(0)) or clr_endrbyte_wire);
	wire_end_rbyte_reg_sclr <= (clr_endrbyte_wire or addr_overdie);
	process (clkin_wire, reset)
	begin
		if (reset = '1') then end_read_reg <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then end_read_reg <= (((wire_w_lg_rden_wire492w(0) and wire_w_lg_do_read407w(0)) and data_valid_wire) and end_read_byte);
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then ill_write_reg <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then ill_write_reg <= illegal_write_b4out_wire;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then illegal_write_prot_reg <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then illegal_write_prot_reg <= do_write;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then ncs_reg <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then 
			if (ncs_reg_ena_wire = '1') then 
				if (wire_ncs_reg_sclr = '1') then ncs_reg <= '0';
				else ncs_reg <= '1';
				end if;
			end if;
		end if;
	end process;
	wire_ncs_reg_sclr <= (end_operation or addr_overdie_pos);
	wire_ncs_reg_w_lg_q380w(0) <= not ncs_reg;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then read_data_reg(0) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_read_data_reg_ena(0) = '1') then read_data_reg(0) <= wire_read_data_reg_d(0);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then read_data_reg(1) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_read_data_reg_ena(1) = '1') then read_data_reg(1) <= wire_read_data_reg_d(1);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then read_data_reg(2) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_read_data_reg_ena(2) = '1') then read_data_reg(2) <= wire_read_data_reg_d(2);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then read_data_reg(3) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_read_data_reg_ena(3) = '1') then read_data_reg(3) <= wire_read_data_reg_d(3);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then read_data_reg(4) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_read_data_reg_ena(4) = '1') then read_data_reg(4) <= wire_read_data_reg_d(4);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then read_data_reg(5) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_read_data_reg_ena(5) = '1') then read_data_reg(5) <= wire_read_data_reg_d(5);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then read_data_reg(6) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_read_data_reg_ena(6) = '1') then read_data_reg(6) <= wire_read_data_reg_d(6);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then read_data_reg(7) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_read_data_reg_ena(7) = '1') then read_data_reg(7) <= wire_read_data_reg_d(7);
			end if;
		end if;
	end process;
	wire_read_data_reg_d <= ( read_data_reg_in_wire(7 downto 0));
	loop46 : for i in 0 to 7 generate
		wire_read_data_reg_ena(i) <= wire_w477w(0);
	end generate loop46;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then read_dout_reg(0) <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then 
			if (wire_read_dout_reg_ena(0) = '1') then read_dout_reg(0) <= wire_read_dout_reg_d(0);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then read_dout_reg(1) <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then 
			if (wire_read_dout_reg_ena(1) = '1') then read_dout_reg(1) <= wire_read_dout_reg_d(1);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then read_dout_reg(2) <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then 
			if (wire_read_dout_reg_ena(2) = '1') then read_dout_reg(2) <= wire_read_dout_reg_d(2);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then read_dout_reg(3) <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then 
			if (wire_read_dout_reg_ena(3) = '1') then read_dout_reg(3) <= wire_read_dout_reg_d(3);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then read_dout_reg(4) <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then 
			if (wire_read_dout_reg_ena(4) = '1') then read_dout_reg(4) <= wire_read_dout_reg_d(4);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then read_dout_reg(5) <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then 
			if (wire_read_dout_reg_ena(5) = '1') then read_dout_reg(5) <= wire_read_dout_reg_d(5);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then read_dout_reg(6) <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then 
			if (wire_read_dout_reg_ena(6) = '1') then read_dout_reg(6) <= wire_read_dout_reg_d(6);
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then read_dout_reg(7) <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then 
			if (wire_read_dout_reg_ena(7) = '1') then read_dout_reg(7) <= wire_read_dout_reg_d(7);
			end if;
		end if;
	end process;
	wire_read_dout_reg_d <= ( read_dout_reg(6 downto 0) & wire_w_lg_data0out_wire446w);
	loop47 : for i in 0 to 7 generate
		wire_read_dout_reg_ena(i) <= wire_w_lg_w_lg_stage4_wire443w444w(0);
	end generate loop47;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then read_reg <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_read_reg_ena = '1') then 
				if (clr_read_wire = '1') then read_reg <= '0';
				else read_reg <= read;
				end if;
			end if;
		end if;
	end process;
	wire_read_reg_ena <= ((wire_w_lg_busy_wire1w(0) and rden_wire) or clr_read_wire);
	process (clkin_wire, reset)
	begin
		if (reset = '1') then shift_op_reg <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then shift_op_reg <= wire_stage_cntr_w_lg_w_lg_w_q_range103w104w105w(0);
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then stage2_reg <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then stage2_reg <= wire_stage_cntr_w_lg_w_lg_w_q_range103w104w105w(0);
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then stage3_dly_reg <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then stage3_dly_reg <= wire_stage_cntr_w_lg_w_q_range103w106w(0);
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then stage3_reg <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then stage3_reg <= wire_stage_cntr_w_lg_w_q_range103w106w(0);
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then stage4_reg <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then stage4_reg <= wire_stage_cntr_w_lg_w_q_range103w108w(0);
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then start_wrpoll_reg <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_start_wrpoll_reg_ena = '1') then 
				if (clr_write_wire = '1') then start_wrpoll_reg <= '0';
				else start_wrpoll_reg <= wire_stage_cntr_w_lg_w_q_range103w106w(0);
				end if;
			end if;
		end if;
	end process;
	wire_start_wrpoll_reg_ena <= (((do_write_rstat and do_polling) and end_one_cycle) or clr_write_wire);
	process (clkin_wire, reset)
	begin
		if (reset = '1') then start_wrpoll_reg2 <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
				if (clr_write_wire = '1') then start_wrpoll_reg2 <= '0';
				else start_wrpoll_reg2 <= start_wrpoll_reg;
				end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then statreg_int(0) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_statreg_int_ena(0) = '1') then 
				if (clr_rstat_wire = '1') then statreg_int(0) <= '0';
				else statreg_int(0) <= wire_statreg_int_d(0);
				end if;
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then statreg_int(1) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_statreg_int_ena(1) = '1') then 
				if (clr_rstat_wire = '1') then statreg_int(1) <= '0';
				else statreg_int(1) <= wire_statreg_int_d(1);
				end if;
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then statreg_int(2) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_statreg_int_ena(2) = '1') then 
				if (clr_rstat_wire = '1') then statreg_int(2) <= '0';
				else statreg_int(2) <= wire_statreg_int_d(2);
				end if;
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then statreg_int(3) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_statreg_int_ena(3) = '1') then 
				if (clr_rstat_wire = '1') then statreg_int(3) <= '0';
				else statreg_int(3) <= wire_statreg_int_d(3);
				end if;
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then statreg_int(4) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_statreg_int_ena(4) = '1') then 
				if (clr_rstat_wire = '1') then statreg_int(4) <= '0';
				else statreg_int(4) <= wire_statreg_int_d(4);
				end if;
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then statreg_int(5) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_statreg_int_ena(5) = '1') then 
				if (clr_rstat_wire = '1') then statreg_int(5) <= '0';
				else statreg_int(5) <= wire_statreg_int_d(5);
				end if;
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then statreg_int(6) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_statreg_int_ena(6) = '1') then 
				if (clr_rstat_wire = '1') then statreg_int(6) <= '0';
				else statreg_int(6) <= wire_statreg_int_d(6);
				end if;
			end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then statreg_int(7) <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_statreg_int_ena(7) = '1') then 
				if (clr_rstat_wire = '1') then statreg_int(7) <= '0';
				else statreg_int(7) <= wire_statreg_int_d(7);
				end if;
			end if;
		end if;
	end process;
	wire_statreg_int_d <= ( read_dout_reg(7 downto 0));
	loop48 : for i in 0 to 7 generate
		wire_statreg_int_ena(i) <= wire_w_lg_w_lg_w_lg_end_operation502w503w504w(0);
	end generate loop48;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then write_prot_reg <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then 
			if (wire_write_prot_reg_ena = '1') then 
				if (clr_write_wire = '1') then write_prot_reg <= '0';
				else write_prot_reg <= (((wire_w_lg_do_write72w(0) and (not mask_prot_comp_ntb(2))) and (not prot_wire(0))) or be_write_prot);
				end if;
			end if;
		end if;
	end process;
	wire_write_prot_reg_ena <= ((((wire_w_lg_w_lg_w_lg_do_sec_erase532w533w534w(0) and (not wire_wrstage_cntr_q(1))) and wire_wrstage_cntr_q(0)) and end_ophdly) or clr_write_wire);
	process (clkin_wire, reset)
	begin
		if (reset = '1') then write_prot_reg2 <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then write_prot_reg2 <= write_prot_reg;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then write_reg <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
			if (wire_write_reg_ena = '1') then 
				if (clr_write_wire = '1') then write_reg <= '0';
				else write_reg <= write;
				end if;
			end if;
		end if;
	end process;
	wire_write_reg_ena <= ((wire_w_lg_busy_wire1w(0) and wren_wire) or clr_write_wire);
	process (clkin_wire, reset)
	begin
		if (reset = '1') then write_rstat_reg <= '0';
		elsif (clkin_wire = '1' and clkin_wire'event) then 
				if (clr_write_wire = '1') then write_rstat_reg <= '0';
				else write_rstat_reg <= (wire_w530w(0) and (((not wire_wrstage_cntr_q(1)) and wire_wrstage_cntr_w_lg_w_q_range522w523w(0)) or wire_wrstage_cntr_w_lg_w_q_range524w525w(0)));
				end if;
		end if;
	end process;
	process (clkin_wire, reset)
	begin
		if (reset = '1') then wrsdoin_reg <= '0';
		elsif (clkin_wire = '0' and clkin_wire'event) then 
				if (end_operation = '1') then wrsdoin_reg <= '0';
				else wrsdoin_reg <= datain_reg(7);
				end if;
		end if;
	end process;
	wire_mux211_dataout <= end_add_cycle_mux_datab_wire when do_fast_read = '1'  else wire_addbyte_cntr_w_lg_w_q_range158w163w(0);

 end rtl; --altasmi_altasmi_parallel_3kj2
--valid file


library ieee;
use ieee.std_logic_1164.all;

entity altasmi is
	port
	(
		addr		: in std_logic_vector (23 downto 0);
		clkin		: in std_logic ;
		datain		: in std_logic_vector (7 downto 0);
		rden		: in std_logic ;
		read		: in std_logic ;
		reset		: in std_logic ;
		wren		: in std_logic ;
		write		: in std_logic ;
		busy		: out std_logic ;
		data_valid		: out std_logic ;
		dataout		: out std_logic_vector (7 downto 0);
		illegal_write		: out std_logic 
	);
end altasmi;


architecture rtl of altasmi is

	attribute synthesis_clearbox: natural;
	attribute synthesis_clearbox of rtl: architecture is 2;
	attribute clearbox_macroname: string;
	attribute clearbox_macroname of rtl: architecture is "altasmi_parallel";
	attribute clearbox_defparam: string;
	attribute clearbox_defparam of rtl: architecture is "data_width=standard;epcs_type=epcs4;intended_device_family=cyclone iii;lpm_hint=unused;lpm_type=altasmi_parallel;page_size=1;port_bulk_erase=port_unused;port_die_erase=port_unused;port_en4b_addr=port_unused;port_ex4b_addr=port_unused;port_fast_read=port_unused;port_illegal_erase=port_unused;port_illegal_write=port_used;port_rdid_out=port_unused;port_read_address=port_unused;port_read_dummyclk=port_unused;port_read_rdid=port_unused;port_read_sid=port_unused;port_read_status=port_unused;port_sector_erase=port_unused;port_sector_protect=port_unused;port_shift_bytes=port_unused;port_wren=port_used;port_write=port_used;use_asmiblock=on;use_eab=on;write_dummy_clk=0;";
	signal sub_wire0	: std_logic ;
	signal sub_wire1	: std_logic ;
	signal sub_wire2	: std_logic ;
	signal sub_wire3	: std_logic_vector (7 downto 0);



	component altasmi_altasmi_parallel_3kj2
	port (
			illegal_write	: out std_logic ;
			read	: in std_logic ;
			wren	: in std_logic ;
			addr	: in std_logic_vector (23 downto 0);
			busy	: out std_logic ;
			clkin	: in std_logic ;
			data_valid	: out std_logic ;
			datain	: in std_logic_vector (7 downto 0);
			rden	: in std_logic ;
			reset	: in std_logic ;
			write	: in std_logic ;
			dataout	: out std_logic_vector (7 downto 0)
	);
	end component;

begin
	illegal_write    <= sub_wire0;
	busy    <= sub_wire1;
	data_valid    <= sub_wire2;
	dataout    <= sub_wire3(7 downto 0);

	altasmi_altasmi_parallel_3kj2_component : altasmi_altasmi_parallel_3kj2
	port map (
		read => read,
		wren => wren,
		addr => addr,
		clkin => clkin,
		datain => datain,
		rden => rden,
		reset => reset,
		write => write,
		illegal_write => sub_wire0,
		busy => sub_wire1,
		data_valid => sub_wire2,
		dataout => sub_wire3
	);



end rtl;

-- ============================================================
-- cnx file retrieval info
-- ============================================================
-- retrieval info: library: altera_mf altera_mf.altera_mf_components.all
-- retrieval info: private: intended_device_family string "cyclone iii"
-- retrieval info: constant: data_width string "standard"
-- retrieval info: constant: epcs_type string "epcs4"
-- retrieval info: constant: intended_device_family string "cyclone iii"
-- retrieval info: constant: lpm_hint string "unused"
-- retrieval info: constant: lpm_type string "altasmi_parallel"
-- retrieval info: constant: page_size numeric "1"
-- retrieval info: constant: port_bulk_erase string "port_unused"
-- retrieval info: constant: port_die_erase string "port_unused"
-- retrieval info: constant: port_en4b_addr string "port_unused"
-- retrieval info: constant: port_ex4b_addr string "port_unused"
-- retrieval info: constant: port_fast_read string "port_unused"
-- retrieval info: constant: port_illegal_erase string "port_unused"
-- retrieval info: constant: port_illegal_write string "port_used"
-- retrieval info: constant: port_rdid_out string "port_unused"
-- retrieval info: constant: port_read_address string "port_unused"
-- retrieval info: constant: port_read_dummyclk string "port_unused"
-- retrieval info: constant: port_read_rdid string "port_unused"
-- retrieval info: constant: port_read_sid string "port_unused"
-- retrieval info: constant: port_read_status string "port_unused"
-- retrieval info: constant: port_sector_erase string "port_unused"
-- retrieval info: constant: port_sector_protect string "port_unused"
-- retrieval info: constant: port_shift_bytes string "port_unused"
-- retrieval info: constant: port_wren string "port_used"
-- retrieval info: constant: port_write string "port_used"
-- retrieval info: constant: use_asmiblock string "on"
-- retrieval info: constant: use_eab string "on"
-- retrieval info: constant: write_dummy_clk numeric "0"
-- retrieval info: used_port: addr 0 0 24 0 input nodefval "addr[23..0]"
-- retrieval info: connect: @addr 0 0 24 0 addr 0 0 24 0
-- retrieval info: used_port: busy 0 0 0 0 output nodefval "busy"
-- retrieval info: connect: busy 0 0 0 0 @busy 0 0 0 0
-- retrieval info: used_port: clkin 0 0 0 0 input nodefval "clkin"
-- retrieval info: connect: @clkin 0 0 0 0 clkin 0 0 0 0
-- retrieval info: used_port: data_valid 0 0 0 0 output nodefval "data_valid"
-- retrieval info: connect: data_valid 0 0 0 0 @data_valid 0 0 0 0
-- retrieval info: used_port: datain 0 0 8 0 input nodefval "datain[7..0]"
-- retrieval info: connect: @datain 0 0 8 0 datain 0 0 8 0
-- retrieval info: used_port: dataout 0 0 8 0 output nodefval "dataout[7..0]"
-- retrieval info: connect: dataout 0 0 8 0 @dataout 0 0 8 0
-- retrieval info: used_port: illegal_write 0 0 0 0 output nodefval "illegal_write"
-- retrieval info: connect: illegal_write 0 0 0 0 @illegal_write 0 0 0 0
-- retrieval info: used_port: rden 0 0 0 0 input nodefval "rden"
-- retrieval info: connect: @rden 0 0 0 0 rden 0 0 0 0
-- retrieval info: used_port: read 0 0 0 0 input nodefval "read"
-- retrieval info: connect: @read 0 0 0 0 read 0 0 0 0
-- retrieval info: used_port: reset 0 0 0 0 input nodefval "reset"
-- retrieval info: connect: @reset 0 0 0 0 reset 0 0 0 0
-- retrieval info: used_port: wren 0 0 0 0 input nodefval "wren"
-- retrieval info: connect: @wren 0 0 0 0 wren 0 0 0 0
-- retrieval info: used_port: write 0 0 0 0 input nodefval "write"
-- retrieval info: connect: @write 0 0 0 0 write 0 0 0 0
-- retrieval info: gen_file: type_normal altasmi.vhd true false
-- retrieval info: gen_file: type_normal altasmi.qip true false
-- retrieval info: gen_file: type_normal altasmi.bsf true true
-- retrieval info: gen_file: type_normal altasmi_inst.vhd true true
-- retrieval info: gen_file: type_normal altasmi.inc false true
-- retrieval info: gen_file: type_normal altasmi.cmp true true