��/  ��^k*��A��D@7�քW�g̝�G�^�T�|�IVϪ�y�p;�5��p:#�oj#�_�����H�+k�6T���C�-fZA!�0{74L u*a�x�@�9^���Ԓ9K0���tv�p_4.}0(k��y�ɨ��Q� m$�zPY��>�p������W5@2+��XS��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0����Qe��-I3E����(�l�����<r��R7���aF�:�y��{�v�L��$�0������l���;/��e�|^��<<B?���D'�HM
�����a��R�d���`u0���C��V�4ް��ę3��dV�'#�`[�n1�|��HC`����,���B~sO��5��!?�Q��^�#	(H�?x;��>��^��a�PD�~{�F\`�V�b�:�Z�@J�q���$K���UÁ�K
�y �Y�90y�ˇB�V:�P%x?�� +'�ćx�
�d�(�`C� ��C���Pcmq���jLJ�W�ALOIc��,K9k�� �(7������3<���"�'����?h��OahAu�i�MXYm9���W�gA�"_��XxqY��JkG��R� �sw؁�A���5����Z��^s�2<���̏��Y-%�/���޻�s�06�_�V��siD��x�
��h�t��u��:�b�%U{���oU6� /�8x���d��s�i��x��������)�D3{�i3��*m������y#�G��}�UI�*}GI�P���ц��d�ĝ���{�2Ͳ�So��&������s��N�j7->[�Mm�*���_^����j��T�$�L���8 �%��T|�nU�s�/�q��P�3�q�kۨ����� L��ߋ}Y�$��y9B��CzQ�J����|L,'��`���k�$�F��%N�z�G/�-�0��2O�f�/iiS�Ђ�>�2��'$�9��+����#�]:�{N�DG����*1�<�Du���CM������]��TY)h�ן�	���Txq�a-��7-ҥy����Ul~��A�^n=���qߚ�'ZF'�5��'�1F�@M�}�,���gx�{�h��x�C+wa�J�誟�G^�?��V�a�u�LI��%����7dxP��w�FE��3�xQV�2]��I�D �C ���zLݰ���oH���S8��I�%�^�F�t��.�%�ܺ�vU�]]� A�d�C�����.R �})nŸ��v��T��8����k5o��;�{9I�dQ�{�K�|��B��i�r���hA�`?͠F�GM�����h�	F2���� �ze}%��u#�"��$XomP\9�® b0Y7Os%��8�Õ�y�Cwq���_�O��WO��J�8RkЧ૥t��.�ח8�b2��?�="�����1rC>�`1ο�*�<���:��b�w�g�4F�"$�S��|N�i�4T7�,���M���ؼ��5Q���I��
�y�Yn.��� �aj��
/���v��U)t�$�&>)�,��1��J��rZ"i���A��^�{>��Z����%�������
2��t�<���5�u�E⢞I��Ȱ��P�:ןL �-��u�ؾ=�Ig�W�q͗h)�l�5Z�J�G�W�yx)�)����1:����6��E)JZX�+��(��4Liш�7[��lK����p�:��5���_�S�bjZ��ش�JBs{R�6QZ��� �{�����܌3Ogq5�vB=���ڥ甧iD�B�r4a��~�N�g��.���� ����@��~�5�ӓ��� ��|��U��B&
.I����g��,�vd�A5.iz�`���{Gh⡦̴^h-�=ҿ��מ�+�;���7V�E�@H9kO�M�¨5����q���j� `!T��[�rQGt1u11��A}xq�˪��:`����)M��8��B��j�_Щk�n'�l�x�9�Yנ���z3?>�/�AS���Z�T��SsET�p@Y��Xw�Y�"
���Q�4�n\�.�g�6ó+܉���V�Ǜ����L�0�[�.�5+��# #�Z�[%=1�N����M@����I�Ȇ|шb��4���aK�o:�P�
L�](m���.m��)+���0c��3���ur�9<f��k^�#�?����1a}��4*��K2���<��V��z�7�������1y3s���JD�2�S��B���J��^�u�Y���*��S8]��UQ�.������~d�j�>4w4�	�x-�T*��8��U���:�'[�4�T��/~9�����
�U������k�����8���q#N�4LR�撊��*��W���	F�,s����V(ͩ�S�G�I}�@6�������$�ᦰ K�G�k����p�L��!���yɭNz�z�_.�0�7"ܘ�,eǿJ���Dѹer�h2dz�xh��Y��i����Ҧ`�vE*����Wx W�N/�N���H���ǐ��as?M���<���&��ܱ�!s��!��t����$
�@���E��H~%6���3-��]E]1g�<��C��&	�^Gj���ƅ�a�Q�V��Z�8}:D2�0P�׏�%��f��'M��DD���^wX��4�N :���A9�y(o���*`�ٷ�j,	F}� �F��#���e�
'��X���cRfW*\z.���4�p;h�~���������?���w��=j�]~c[�K�i�`�m ��}?���kek^/�>�*�c��K�������|��Ckt���o�/�� ���5����V9�ݧ��=�_�/�bI����D-.������gh�Zfav��d
ғƌ�
)�󕉙k���!���R��s�)W�V��:�Eڔ���Vyp�m��W��.6x� �sz@��M�Jk����"�N.������b�,��p� @�k���W�m9q4)��c���=ϱnE���3{��ڗ<]�c���/�8}0G��$�a~T���v����W�ǐ5���4*�pT�.^�;�T/�aGxAA�HB^���w��}ښE�4�?�3��i%cA�i�袈������ߘ<E�!	�J��О��\�Kݢ QC��K����ٝ�ʫ�S%D�$B�
O@$���`곳�{�71з�Oe��t�����< v�&bĊl;�q����~�����AT�D:?Jr�������>��(bS�6�i���N=�Ivc��xi�h�4���`�r]ؓ�D@�e.�5��� �+�o.4��墾����ڒ��5w�@o�)%8�X�/��������9�,�~��L�ظ�s&B�q��3\��z�Id'����t�o��}��)���*��hbJ��'o������٢��}�[~���q
��M����u��i���5�Jn(ܛ#��z�g�Pz�@  @<S��W�M�R�3��qm�`o�G�Xă�2u���8�b�;�m���@���=د�p��
)���qAj-�i��ɜ��{G���գ��Q��d�R����-8!^ܠp�ݡ��������k�z��4���}etko2n�ڶ�'ZC�!ɥo5�X��=/����&�wP�A��;mqq�	P�:f�E\��Ë���j������1��k�{���I�[C�T���)�J��Q���`�#�w��-
iݖzm�7W���uL�l���mCJ�f�TB�!~♋��c>?(�ca �⍻~7f��1��3���1��պ7ԇ�	-�"�:D�`�9�=,�3l�0uXR~�5/Zp��S��Ze�v��j���s�}ځw�:���Y���ጙm�y��`�%UW��j��<GC�_'W���,�A9��'��`OO��p���Т�(���!h��}�nz��k�pW�� )������,��Ai��O�'���"e�2����;����v*���s�&L9��#��~��!�5_9Ȑ�h^�W�k���E��W�{�{�S׀��g{�����%��$�<��1�?����=�<ی��s��GgID�Ӻ�P�/��/3�P�n�Z���&��*��d��r��2.�;n̛�ן�#��
�C��gg\��n�Ah��X�ڙ��D�jSވ�H���#��,�(+�v�X��*vXb����pX�N�7uEF��>��;K���{:��e�`�e*�����S��Ll|\:���ןzVw��s;<(�:��P
h�#��*�o�pǨ�z�t�k�8��I��
9�'=TԐFhǵ���앩�.8��N��^��-��0����}���\��vΣwTe�y�HNzi�����s��k������>6�u�#���/%{�uy,�� ��ʶ;s|_Π����-�{�����ȟ�������-q�L�U���c��Ll�P����]9�@=A^
��a<���DJ�7��Kx��7w�r�`T��E+�U_�JY��e���z[�ۄ$�rML�ɶ����y~��\���򧔹�̠�S{)%�����G{���Z��Y�:����n%/F[�(|7X;��Z�P�����h��kf��L1�;�ь!Q�A�$�d�0kG�=���9{�})[����<�:�Bq�h4~Ѐ��e6|�phzc��;^Gk�2��MS=!Cn��ۼ�����RP�}�L�B�(X�������˝�C���T��p1h�� �����+���;_��O3㿄�R�W	�%�U�2[�z��0�C�Dw��ti��!e��S�E}X���_!©W�G�V�:���zp��{(��)�"d&b��n��wǻ��e-����O�#�"��k���"wj�o�� ɩ���o��6�3��H�Z$o�c2JsM�z�(�����rۋfB��������i��+1�iO���
�R�b�<�a6O��v%��al�(:m�~o�$؂1$�0��/Y��#
�C5���'�f�O%���A�F� ��_�Rއ9�񌿒�}�J��bu�vc��b��C�T�&>Mj�*���^fL��~�t������W���kn3(����,j�M)�/�o�%4�G/ա��T�iR��v���_j���RZ��_�7�S/z��[]5dݢ0=n�ǅ�aVj�Lj#&�� ��n`tY�V=մ%�$榧C}�Fk�nx�ot�z;�tl���G����G.r(�Lu�����o��s�۰;�G7>Ne ��~�A�ooO�|9S�LpzO���d�s����)��]�j��i&���,a��a1$[���2��M�#�¶�E��0��.K�L:�t�@E�P�=��O�V+1���< %�i�{����&#����ks}G�[(Y'�<[q�w`Qe���ɈH�$��y�W�=�նC*��Ҭ#�}G��UG~�m>S/���{����F���pI ���#��1���[(i�3\�9�~EWV@��`4�:��@�����!�40����E�8�/��kYU�I��6����G���u�\(�I��	���1<�QL�B$�^g�V��mC�s�,���[ݒ�cs�jԹ�po@�1��>m��8��	=dX�c-�T'R��M+!�p=3o5�'e#�Cԑrc.�H���vV�;�u��a� C�*D4ɑ&�P����綦�m4<��K�ש0���5+��)�w��}b��&X۬�n ]����9o��vZ��д'iGJ?(H�u*�~����V�S��A�Hwtg��_�m�)8 .�`���7���)/cݢ�Z����>6����T cu���"o9$ ����Y����S̈́@r}/����
��ߒ���:}(�)cC�XF�I��G1C6��E=��F
��,����}��,�g����
r�4j��??>Z ��{޺���vJ�\�����L/�z:������P5Y�	���K U��4�&_��Sx�6U�� {r�#@EF���FWtC��� �:׊2�.L�^t�ʤ��A�6���5�"���W3�����M	Ŕ��?q�r�YBJjy��$���Zq��}����cʃ��}�F���b��rA���yyr&|�8�\X_*X+6��Up��\�`!�����CJ���
�?Ϧ�s�F�4}J �]E�JsU�^�9��#�w�.�}t�m�xWȇ+�r��t�t�q��f%㺽��:u}�cM�rX�jgi���^&H���N��&$�OV��X�$�����rn�%��ѹ��J0mT0�$���0��3>�`$�i��F�����$��u���;�֖���^���z�0	 � ��VA',*��v�W�˃z�j*��_a����#ЋU�/X����~7k]��,���b���+�e�c�&���l�נ)����LǛp/�$�:Dm�g7-Ǽ��2Pb%m{S�����}6���a<�%1H���g�2E��t[��@�Y�����N�6��qT,	nx�|��L�ew8�b9	����o��.�=�Կ�)@P�רz D1�,K
+ ��i��x��r�b9���2 T~�gms��7���'�.\g.�6%��q���C8k7ڌm>��%^�ٿi��U!��߿ȳ��w���S�� �q���y��3h��[�+�y� ��� �����_� ]�?�)8��oME�	��v��jt��q��6�$4dU��B{z�}�/�7�`��T�@>���
r���7��A��* 5#�z��3�,V���a]��#q^�� 7+	�����UVga=�x�ٖb빢����j<j��*���´�;�շ���+H����\�1��+�*���&P�ۼK�D���S7O�s�+L?�|��= ����0��!�7�*Ar&�+�Ī��ǧ;�tH'nr���K�������UE���\�Z�őAm�����(�n�7u��xl Z?>�i�:th��G���?���/�QB��O��5��K�5s�&�;S=s��e��:�W���QL�{h��nqq��!�p��D�����IƏ0#.�GWv���D��aI߱ӥE�{ռ�b�5t]wE��r�������:��:��4����Y	��|��ZP�AKK:�̴@��[b��$u+k�?�+��H|�p!�n#��iS�t�����:;7�-+���U�T����h��?u���;��#�R�H�Z�v-2q�����f�� V^�����g'��tA��� N�2��q����0S�����ӠW��)�U���b���?㪝�7�|ہ�F;zm��C�f�A�0�v�'���4bB��Xԫ�c���ܜ��1�vM
$��\%�]8��I�~���T����������o�bn3B�������=b/nf,ŰK�D����ښӽo������Ԭ��4���7͞�~�+�?�#��l�&�Ii�V���p�3.4��[ݷ��Ǵ�<W��$m5�W���|�Q�Aս!���X�'��wθQ���Ջ�F�1�,��$jo��a��g��������8R�-��'�������9�e	l�vS�g��6'������C����V�{���6���WN��A4���$%�C33��<c���?��.����/I[S�y�yu]�r�-x�`�����%+9��5����)%TK�5��-��������mL�4$w{��%����` ��hz7�S��3��4=��P�J�T4�eM�r��8�ֿ���'/��HI �FL�	��j���JjF�V U�+b*�)=.�L%�`�f�?�S,��᷋,z+��dhUE�ߣ��0���Ȳ�	q�\\XN�M�̬��x5\�&���Qw^�=�����'O��G���\j�Ic<o��#w�[�Ŗ���G�8�,[wy2�܉�B�##��ʄ=�ø���u��p m�zؖ=[�oW�|�ī�~��,|=A�TZ����MÒ#�����2�,���YQN݌��J���}�`����<4��v��֊$<h%K5��Rs�w�)s�!r�ߤ�j^���菗\�-��2ܔ{�S�?���7��Ysa�Ժ���iy0���`��M����_�S�2�>*��^�3�k��V\Pl�!�O;;f&Յ�+o?7i�͇7/"ڽ�h���i�0C[P��(0n3�V�=�p~=�[�ąj|��"$��+�~�UT謋Pch�ɜ/A����ͭf|<�
�)�X�4�Rn(���U��\����I�W9��`�E��jt$�k'^���`-�7�y̶Kı�ߕ�:m����).JT�"���6'-lp�#����m��o��:A#M�!՚�3"	"e� �I~,����y/m z~h��������yh6(V1�d.>�CE��(}0B�ٯ���r�F�ft4t�~@�l�b����r.9 h���,QI2DЖ�k�&�	BXӡ��|!a�"S*[���<��?5:-m�H�~F����#�/�l��T+F�70r��Ӹ�����Tce��d8A4��u��}K�<�<.AEa8��RVK�!��n���Ec�y�D�&fNs������U���P�_�axY��`��3�s^���|���2��oB��G|�%�dZ�q<R�拼&�����R���Z&�l'�
T��:�D�Y�B,ъ�e.�����Xex�g>�Nİҽ&׎>2]SvI����?茟EE�٤r_�'K�����fD	�@���c�Ӛ��3�����:~���zp�	et��AW�q�.�O�#|�y �h|h��u�h Ǝ0�4|�O�g�+l��E��.P(����}��� ��Z'�J�D��%6 �荋��l����xN�������RH�a	g MXxO8pn���	��C� q�#5�%	�%ka�ބ4�J"!]R�'�xN��7��_0��B����LqWپ�y�hK)�(��o���U$�W�-�~{���ݠ�Y�^�H���K ]+�۝��u� ����M�Y�L��ZGz�.����&A ��1��F�dy�� �!�Mf0��Da�H��I"��TjoO$у��A�����'� Ю�܎�rk�~���#?[,�y��L�8Z~��&��"�x5���Z%>��t��#\�zqO(
׷me��ܝ}8����Iک$��70���8��do_�=Ӷ>���l�_�}z�M�y�G�^8
r�Ѧ�cK|S�Q(>dX��3yc9��r8+Y0���X�C�c,+�Pp�;����B�<��P����Ҋ�B�߆�*��&Jm�p7��f;X]�#4�DY�X�6��b��!^3��RP�:�rF�8��,�Cͣ4|��dl�4���O� ���ڰ������0�]��ة˓w���������4��^" ��C]��vڼd㈽_"AFI��u�
���e�C�\[sY�:��>�i�>�w��������א}��N��m�������n͓��h�q�o��9W��Ш$aԘb����1��L��h[��Iy���h�Ub��x/.ܝ�a�T���"AHm���s�X���m�/�>�XZ���4�LP�sK�W�� ��(-�U�;�|�֙V�l��eE�D��[Y��))�����#���O� DJ��(�`H��ӹB3D�X5�-}��'��+�3���>�؁��R�N�k���8���P!�u3 �;5�^��U�qQCMp;W��'��3������L&্�d�^�L��T�a�
�(7���5+���߂�&��Xs��Q�M������$��$F�E�*ݦ5�n�	��vϵ}#Od��^̤��Y�m<T�����+H�����d�B� |��|�Ț��A�,M����s�]7���]�z���LAQ�GHͺ�(�[?��������с7��ޗ�N5��@�L���#��Qf���$(����į���&3�U3D��ƪ�Sg�~���fh�.�"=��W���DN���*�K_�U�z�~��Z��)}�ȹf�Ǆ�'�aB}��ɳkep��!���쫋0y�Ӧ�aT拑}��U��i!J��Bz�Ē�A&�e�U%Ng#5�o�����]�E\e(=2%��L��\ߧ��ρ>�?���V�m�R���o�=��'�9�a�Ƕ�� fǒ����_�~��E�����R��z�嘪�%8���C^��0��ز.���أ�{}f�a���ǣm�Ė�q�oZ"�����_g����0��Uu���NsL�e�)Ӂ�����p�.��p��� �\�Q�B�z?��ynqPe��+]���!h��= �9IM��)r��N�_�um�%ב.>��{�d��k�{��]����s4D����YndH�p�@��lr�������M_��	��c����w��|KԘkrP��ޤ�G���e�m+�
H�]�����nm�
��Р��5T9��CL��u�Uh����H۷����f*k�����:��a�3�=��½'n��^.�^f"�/�τjP5%�J�~��Ch^BTBU��M��w^*R�6���m�Ո�c=��t�3�3��u�~��q'_�*x�b�5Iۉ�����\({��>/�h�}m��K���k��ojJ�٥m)��n*�Sq+�#���7Y�F�.g�Y-�h+�\ʟh�0`ku��f�Gl���
��� W�dla���%b�j�_�k���gl�����m�3�
�b��R�`��L��ҧ�v�PÐ$ �ص<7f90�Rs+���Y�T�T�ͽ��c�2/m��@���@���;q{��h=)��&)t�2�D��E����5@W�c�P̪�ݾ�)K#�p L��	��?B���M������[�C�(�zLu�#6F->�2|d&m���8J|4PvTJ����k&�Ol|�`%	�
��#C���%���]�aC�Z�t�)@'@���=`6^Q�D�]���`�/(�+T#�D��o��G8���.��ls����g��n�|����}&i�dJz��&���y(�^��W�iK��N����)�XKHʲͿ�* &;v�����&�4"VM�c�>�"s���h��A-�'8�>~cC�����W	|��+�evNP��~����W�-�/a��/���/�B7�,?��r�>TE[���N�@h�0
�|�P^+�����(HjgJ�̀����VV���n��b�d��JT;M~��gJHKq~�0M2l�96:9Jhi��r�LD8\���!�ykoT=tp^�J67'�s�4B��Qtb�)�b�5z�Q��:��_H�@5C���+X�9�<}�9*>~;^�M[R�c�cD�[�M�S�u����_'��������N���jz��$���8wm���qFD�E�{is����gB�p}X������E��?.G%�D�9@�kq�Q�#R���4g&e|�}���`��6!~��(��(��%�ѐf�h�"a7�J���g+ӝ$��QTo�D�s��}��f��,H����尟y��h��<���aa�Tq�b9�������J�K5>��>&-0�=Φ��":�B����;��A����V7�����h?jK �R�KU�q�L���d���?ֳ�9أ�0I)�k�FvFӶM�J}0�VHB�N�M���@���(��0JV��?�OZ�ũ����J�u$w��l��:�b�yȌ�3���5�B�rw �f�э2�.dC?}Bm!�"4hީ�8A}3=0՝>����-Z	Q򟈲�y�̈�8y\K�'�C��C|�hɢu-�UKa`B��qr��	N^�BnH����y��$��c� 
xI����)ۇoަ��SU[-���_�;J��f�#"�1Ϧn�}	��}A��7����6��Y��>\�|_b�u�G�d&`#���1�?)�J\Q2~1	I��ϖ��vޱ�.c��S���������8B�!��g1e�2TqJ��4ţ��O�$6�Xu��n(����ܰʃ%f�V����z�,൑i�����rv��3���q�Ӡ[�C|��N['�g�ZH���<��	@gX��R��q�0>)��#�	����պ7���;ٔ}�2ZۛX�����{`9��IS���3�w��a�����=��� ޲�DsϜS���c)��I@~Oo�+5����Z6��]W����Z�Δr[W,�H"O��G8���u����e�`�h,��EQ;o�\��{H�r!�I������9Vi�����)��1jkv�a�aν���ȑkr
�.P!���d�`�d8&ظ��yOC(�~ffj�����Fl�;@����>>��4_�q�MU�^�ڗ���
?���[X�U��̝ :�W�!�w�KZ���5����3 {9e�?Es�\�z�3��P�5��0�K��,{�"��iu#���E���q�"��ie�0�K#?r��r��&�ϧg�cS��Ʀ����":Nf��\������Ϩ��,���RD;�k�SU�k���x����>��͡���)���q���QU�s�^�<�<i؞v1EOz?fR��]^m�#Z�0��k�6vE����zˊ���`�o���	�f�ą�/����St|�wT��X�bqzX)�A	_����6�dOI�ɰ�TL;F�A2����z�g�lk�I��U2Q�#W[D�QZ$� ʊ����all�*#����Ty6B�ߝ�k�G�����I����!��'�A%���\o�&{�L���L-B�G��n�����z�t�\\AC�����prD���,$�������7}r�ޙ�O�$�W�x(�z�7_%#�����֞��4��,�T@��?�X-t����Z��GzÁ�t�K��?���^v*4�Vd�� <��#t�9����la��'���%[�c9��vP��r:���F?���	,����(��J����>	�)km����p��@A���y�9ot)n��c�iW�"dIbR��d�����e*q&T>���?8�oܲ��W�t7>Ȼ<��ꬳ(KK��ԡ�+xC"������^x��YL�r\G"���
2�s��W�hsu���΄D�[�Ү��Rj0�3��Ƶ3�H�+��ȏ��K;��3f2��v}dQ�1�M����]K��,*��gRnnSH%��H���+,#���<ߍ���������	g3�LL���!R�`o,�<
���X� a��QӃc�v�&����6SW��dc��Cn�w�{�h�Z!����7������;nNЍ���=j8��*5th�20]��X�W�
V��qJɺ\D�	kt�d�,ߜ������l{�Lm\ɗW��� |���v���|���|��t�;���Qbm���đY��oE�c�հ�i��ͺsY���.nR��	߇eXfZʑc�^��R��I]�����2x|�_--�����+�@�*_��Qj�����U��r��Ic)��C?�୨���݋�Y��e�PWA	�8�
o�6��UC���lw��ʜ�MM�H_�1=}�$���d)T�&j pw9��
B}y ��ڴ0b�D^�Dh|�fj$]��Ө����'�.����`��`�+E�ب�&]��Z�����a�0��
Kz�i�hkE� Kr5?a�PBp��l��l��9�Y�x<�ܨ�ѭ\S"{w�p��l�Bwn-��!S>���kHG�0휺}|۶�<��	�ړ{?S��cnEiy�����%�E�Cx�ńm.=ѯG��Y�F��G��Qf��w�(�J���`������}>�Ǿ}���������O�
i�FY�woAc�y����,�sSb9a�#'��LȺЊoQnb3��ki�:�}Ob/:�(��<�n�3�9��p����a	�|��@�{+��D�����ȏ絊vP{Q!��;��
}H��;Xή�3l$�������AЃ}�����@�Ő�6	뿞�n���b���\��6�*�l*/F�E��[��X�'����4��G��Iǃ�
�' ��
͙����v/.4�?��c�/N����sŵwƐ<���E�Z��y�y��J�h��>jT�?��y��* kE���j�V�(�An��Љ�4�Q'%����-���9:4Z�d
�p����.����Dg�2b*H��FF|A�=PS�m���I��#S^�!�cI�[���"9U[Vu�͹Z����Je)��VD��A[�v�.<����rQ����[�ǦC�V�#`f�eҍ�n��\x�2���E���M��'D���ٛ�V��8M�'��+p.��kAo*�����A� 	���^7�+oXb@B�Ϳ���WL����9U�p�S�����~�O������كo�t<Ѱ�)�����kC.:�a�e5�1O;�H���&� ���Ϩ,�)*��� ��蘞��j�O�@5��P�3)_d��G�}A�q6�)��x\;_��%��b�VG>��փ��x�cu��G8�8q�*����5�1�n AF�;�hPP����%�8��~�Q"5�<�"Љ�D_d̴�k������aMT��PN�D����a�b#De�<S�����_�u�=3���"X���pcg��гW	L4GX� h��?&�)>��&�{�_�X�1��׀ҥ�Ž�����+!��Cޓ}����un���b��^�1~�`Ȍ�6�n���f\�U�M��(��bl�)`�0��)�����)�x��o��YS��9���	��Z�0�1�5����Fx�_)�����|��A����$����*��k[�>B�m�+,d�z��5x <i]��H׭T�H =�%���A� E\�b{��d�}�O�����:"įx�rp.{J�������J:�%B�s"��{\�~ϫy�~�ꘚ��R� ;�"٠�G#r縢��כ��A�
6�CN��ha�Q���^�t=�m����T.bZ�� _�#�]|�;}���Ds�ˠ��_���)UK������ 5(�������r6Jb	��_:�t��Xl�ib�>���㋔{��^����L���6�*z��=�C�+>���䛒��S��~9��%L����GZɠ��*n��i��h����_��k�A	�L|��H�z�h��l|�B:3��=s��V��ʼ4�~���(�b���'n���x��/�2_<V҂�o���BRa��i�T��*��Svu$U���s�b௎�A�X�R�݆u��癑V�b1Y{��AWzh#-1�� ԣ�wB��c�����K23��<�/[J�3����8�'��e�>O�Դ�w���A�/\���ܻM@���������!�B��%�h�c'd��X0�+�\ή�W&�(?=V/�㾺���(H,Ö���Z�Z
W�'$��-"b<'�FC?f=����H�Uc�@���l�W^Hhѿ�}	�x�tk��E��o5F��/	~�BP�#2�q?��}WǮ���!]Zf��;d.��G��:�p�I<E>��H�['�w�A��f�7k����������hZ�B���*�>�v�4�Z��.���.�p�(�گ1C�zJ�1fY,=��M�
��w�+���%]��w/<X�
jt�91�9�t#���Kș@��F���K����z^D�ӗ�r�#�W�P������Μ�ЄI��ծ�.GZ<D��f�ٜ���aV���M$������L���51��s��֐�@�h�=���gǻ@�Aϔ4l��3T�kh��u�g��i'<�w��\�k�tPl�#R��.S5�;Z��4�͉�9�k���k׼�
�=:U"�����^�F)!��	yt�q`��E��#�h`�����:��a�yNv/]L6��lc�V��Jƺ�N� 7~�o2�o`�����@#��}!i,]����:��=Hå�+���H`��&�G�X�V�3�Va@�f� C	���R��V�SHD�2�
��у*N��LNG�R�����1/���m���{�`��ȃ��u9-�i�7���\2��^!|�j����`�<ߩa�S�I?J1�iǲ�Fl�V��Om�w�r� �E��YB=�I��9-�C1�#/�#~Ե����Î�Q��8'��VG ����ɪ�M���[�H�BL��ӏH�W6���Q�!���d��S ��S���z�ٜG��ޫ�j&�7z�?$�2=�<���Ω�v�;��@α���Ơ�n������Y��� ��Vp=��
[�.�ݑ����������[�͕`<�8�7}���㮬b1������W�q��Z�K!�ј�y1� & E�5B@?EF����$GD������nĹ*X�s���ab��|��7��l�U%r��Q��D�?��w�T9�ј|>%48~�z��b��#P���R�g|=4�wc���7S �i.ZN�/:)U���Yɬ�S���i^�gT y��gԝ�e��=K�;1r�Y��jD:Fg��"�x�$�E��CP6��Y���ܪ1�������"cY>JWy1VOD)�Ex-��,���ي��ׄF�U�a��2��ָs�����'Jd(+	:��f���f)��2�)�iL�gx&\�k�9�t8xa�����~��M�5J����9�m� �)�v���I�c�e#��B���x1+g���MO2ڷ�q簏ەh�ǒ��]ţR,,�y?$g)���QGSMF:��2D�\�-s���k����O�����z��0�6�����K����(&o�B�S�t��`�i�y�jt%4蝨=y<�@_㳫��	���~N��;��S��+�WX}S%���vFGGs6
���/Q����k���2&׿���.�e4EV���=d�{�-��ڠ!#Dn`�R�Ń���8�C�}��,^��lF�?}s���Z�G�Q�̿��XL���	���y[4>�{���#�T��#9�H�8P͒�i ��Sb���Dz7�� R�h<}��Nz��6�.�[91my��h_������\QVC����R>��1-e�)
��2l}�|0�S���a��|�i�I��۶ѫ��|�+�������T�8�X?T��֫�46�e�:Uicp������-qޟ��o;*�l(�hi��:3��%T'4�Q�MieGb�YZ&�֜���%O��[���������+�im��	������"�k�7/ �uc�4��]��V����F�.��Nћ�c����ڙ�se�ߛ[���03��f�?�V��`�����q�&�K!߈��	�-�:�,mXȥ���7p���8�g?g����qW�O��F�;ع<F�Dg��p��$R[��S�?n2�㪋�M���?]X���P��#]>��zq�G��Q5�H�m�mTѠ��H�������0X �.$�0*o�a�,Of;)�R5)�θ�}&����*__��S��������ת��:��7�<ү=�y#��[1����� ��+ϙMg�Q�>yB�6�灐/�~��J�]Ӡ�y�%"�t�xg>{ʝ�g�b@K8����6�Y@�]D�*�
*�	�"���n/(��<�g���(oJ��x��$��-f�@�J�q�u&�pU��բ�pq�vؙ�(�j/��tay���P�7=���3�I1Mƭf��TE�Z��YyX�0��r�%`L%�~��p(�#��*�D�L�/��Z�F�.�Ce-Γ�������P*��s�X����i+��Zz�rR��s�������N��E��ne!juN�o}��W����;���V��"!������"����� -� �ߠ��g����jA����$�.�铝7`�5B���D-��T��&��:��!���`��U�WFot�5�*l6����c���ݍ��X?��{�l_#-�a�B���>�٢�s��JF��R9bzV�u![����?��L%-�zkk&�1 �_�Q��~��=���f����0b����y�-�� ��0���m}�y���x�����=���O=��/29z�f����s?��o�q��ɯf~1/Q�x!&������A����f�o8�R�L�F^�W�T�͖��: �ui�22�K�h,JT<�z��;']n������#�۽������״1�{,�bϷ���\�%;��tDEN�s��-'�9�P���_tѮ������d��qf0����@�֞n���n��?��k�;��1|��!��ø��iu�y��t��!:m�WՕc�;C.n3�!�Q]㨗�����������刀EcQ�#��ŸQ�J�B]Ջ�Vٲ� 3=�S���{�/c�|�8�P������R�X�Я�ؽ��ԁ�Y��i^�D�)��l8*�_g����w>�-}�����oI�j%����zT�.��/�!�L���_8����1�v6gnV�j��Cxv�_`����Q���c�sˆ�&���]G�g�Lhk��Ax�#��B�A���@��T@ժ�=G,��X�bC�UH��?��˙��g}n��ţZD�T�$�v_m�KС���cA�V
��Y�6k��/1�$	�'S���Ҩ���l�a]T��G"�a,��)ry����I�n��G+�|�S2��v�� ���PJ� �W���(H�3>=�Յt>�ܵ �'h�/p�EEK�P$��`��I����'@-2��9�Ϻ��)�#]vQj�O�*���z�D��Fw���|�c�E>���*�7ў&Ol�W������ո:>Z���iOK���!�7�0���[�jj�����-�ҦL�%��	9��8�{!5�F��ls��Cg��E�N�Ly�ܘ�M��!�л�^O*]�9g�w���]�5j9��-����D*1Z���]]����+��~^�L�ȝV�AT�8�n��u��5�v����p
&f����;G�+���mc��z�C0���(ܭ����m X���`u��-�׸�Ⲭ��Z%�z]�v��ۛi"�%�8���$*����+6.c�2����Q<�oU�lK�U`Wp(0 	��I�p0m�8��΄��I������q��8~Xț�0Hɹ�B	���;�0�"!���%7`M,q��g@ʕBʈ�8߆�uk;����~>�$��c��� 9%��͸�j�η�T���l�
1�7�7���7���N��v��$��I<A� �^X����&�s��Y�}y!����{oH$˘DN��˛Hpz��o&��J�T?O�i{ko�N�v�3/I����G���t_��A���]���F���l`�����m��]?��o�0 ^l�è/�L�+�幘�+[���5����(zv�Qs3=��UCP��D�T��wܾJ5:�~��LJܑ�N(l�\����W�2k��
����NA�?���1';�Y,&oVP��%LԼ?�q��j��>��<��5Ӏ.E��B\��ܺ,E���J�$v�Q�:�o���c,�[>s�/�-qدZ�7���y\�RwS�.�kaM�eq
�*����"�t:�!�f�~�n��_�Y��"6R�܏B��e5���PH�A���.��\@�1l�d�B��s��(EF���J�%�/Uzw.V�[{.����H
�ɲW�n����DΈЊ_�Մg�%�i���\iG��Cu�H2��K�&�h�mh���V)�Eh�T�!�E*fH�	��K�]jף5k�2z�k�$@���O~�FE4훑n���b�>m�Ų!	�"�f�؄I\Z��IX<_���P�=q�T��ȕ���D��N��R��c�JV��Z#�ه�t ��~M-��5�Z���49rs��;ێ��X��AT1R�p{|l���7���4����KrU"�o�T0���	�.i#m�`.��^B���D�R�8�Zݪ�N�I�jð�y̈���5�����%����������*�Ut.����4	�3��l���s�V���U�~�kB+�]{��A�20�?��=XK�b��y�g��Jg��ұ���	�mÛ�Ϩט���D����>�}�.Ï��h����JI�G��1n9�!٘�<ȈaR�S�*5��\n�/�r�	��d�H���;�<'k3�{�5��%���_�(����u�&"`N&�
{륈�yBiP���T�h�t7���
X�dG #j�qx���v��"��+�W�@v|�FfVa�J^Q5�Zk�w��
N'�Mt�#�-�LqLI:l5A�*Hq�G�����<�X�;�y�V��i�F(�l�B| �S��7_Q��������y�����;�D�Ư�;�"R�k�B '��F���`1ܾ#)s\�O�m�\+�9n��(�2m�a��gA�x�^���	���$���3���h�P*Fv�"��3D���?�p�P���i�q���e:�~����?ʣN9H���X�r�Y�^��3�S���dW�rI� �*৯���*���t�7r�E�l �>����9�tњ!\�]E�	#\�Z�c���j+�4���<�r(ٗ2���H���g��g��\�Wc`�ٱp����0.�傹�_���$ͪ��
`r��,�}�pGŪ�2���rװ���c���y���]�=�ZXDr�W�Boz���]{P�)��}���f��`Kcb����~o��XeӲ�վ�Ymب�$aN���E�ls�|�����`�U�(Þ�Kz�V��
ƥm
d�|G櫞 �V�-�����I��$�Ir�x����R$t&�B!���\�H�Pf��VUv�N4A���E���G	]����"#���k�@6��i���<��R�.��
|���4�ϑ	����YS��$�:��0W}lo\��X]Ek�E��CO~������-���QJ�-��[�r��6:���)��g��F�mH� `֞~�����l�t֪S��_`���~9gyeS� ]��xx�6Ob���yT�vթ��~aT~z:���ڶ	��4;M���_�� ��=-0`��>bO^K�ZX�K o)=�"=vM��.\Z�G����a�7C'{鍁#+�#k�]������&$��}�F�Q58z���K�G8nh:F�)��l�w�N���������MB��CUz;u0�a�
�t��1zrH��-��Z�3��)���oj2MF�~1��7m�Y>Vh�s��<}��L�5Ҩz�<�MT��0�䑪Ӯ�zkJR�P�W���8�xH���JHTz�GV<�ҵ���G�@)?M{���k��:"Q|9K��TP��`OZϽU;�����PlL+���<��-���ԟi��w�7�"C���|&<v��Ki� �0�ӎ~=8	�Q;����K�$-�Ⱦ�=�b�ЍW�y���OHX�'�SL���r&	�	�H#U��m�k'�l��e���>��٨�(+ww����i��k4���\���ȹ��L���k ��΃��8�a�4-���)��~CCڟ����j�}D�+��@����Ne����mҋ)w^{���3x��Q{	���O� o��0m{=��V�ɏ2A[0
)�Xh힭ϪcQ��1t�-��I�a�l�D<)̒3�)l���:$���B��bT��Jd�߱�|B����DNd���&TFX\��`���sBř���г���D��
2%��#���w��@�YH� �{ �K,R��Zf���.'�O����X�����\ϣ����x�.�C%fF�ؓ����($ل�b��"��~��y�#a3��b�X�h	�U\�/�=unC�jؼ�7C?{����<����b�u]o߼:!@���ɵ�v�@�2�,�+u0�uLar;��i�/hr��$ɼ���'R�r$|_GP�G۶
z��]+| U�'g���zXr�뮲J�$G�������h��t�$?g�3ƹ%�%�����!H �YV�X�����PN����WoK�@ֿYq���P}f2ZG�*���x���x[�2�`]�T]�Z�>���߻m�}���}ű핹k�S��W���X��bF���Q/&r9I
���s)a�[�i~���t/0�N$�M�,�Ģ̇��'�ә�a�Y,z�x�ZC��a��\10�����^9XI.1��m��^B�Q����\���R�q�9�F4��b��䣹w|�8v��n��p�k,�53���G��苯��Ǣ��u�ɇ���_�g�4����蹂 ��BC��nMl֓s��ĳ7�K�P���ر����B�k���wGcf��\'��z��!޷5��h�C����LM$w����e��[ai�i(��*��G2ω�(LE�M��#r��v���eC������l���ESl,��ana\���_�oN�-l&0�w��A���c�[2``�a�jw�����.�U�����g�s o_=֑�b�����"0/���E�ʸ�,���v��d���>w��f�Om�C��ԯg�I�^.X�����u�L���;sH����u�>ѝ�Bt�q���9#��i�������i����ڇED���\�}�rќ�)������V��z�o���.Jǐ�p�G7���y�G�j͇�#mي�Z�T�{�� V���d�8��d�@��߰ڮqc7io�����_��g����'s!��М/��:�dI���FI(bN��h�5hP~��ɭ8�
�x�����O���ec2�6��KŚ�b���V��w.`�Ȝ��{-�+�_;HES�C�۳���9a�Y���m�w(���W�QA�9��3��Y1��\�G�Y���;�Ǯ���G}����M�t�uc�'�8�z�g[1NJ/�)/ˈ�{��]|�.�1Au5�֏19���b��u��!&[M~|�����ӊ0��iE`��H��M[��=�q�L�֜m#�7î
��sr����;Ģ����K��1^���k�4]"�h�z��E2&�1�%p6�!�]I��9_b���3^��|0��55�H �f��!4�E�
�se�HVϗf��͑^�oFX?��d�.��j���У=�?�UBHx[nJz�v�Q�6)K`�;�Һ}�S���4LJ�]�]��Ժs�#:�a�Ůx&sl:�k�ay"鬱r�^1'�6m^�c��AD��`����MjSP��|�}���B���ʏ�������N6p?G���y%n}lN�4`(qb��m�-����5(�*C"���IqZHY�O54ze�	tү� �`�tj���(*a�q���mIx>[0�@�/���'Q0?��i��pmVw.h1XӱyvbF൵a��Ws��gS�'�ӷ�G b��QO���)���~�4���Q�O���3N����i����w"~R�����rc�|ېoK�u�	���-�W�b��:LJJI�/�v��T�Gţ )N�]'��%k��S5P��#f�K��@�}�|*���ģ��������0����������?q��{c�Х���33�o��:�wu�|4GY�2�v KUM��/��L<�q�3Fd$����n��vS�]��+��]�z]R$���x��m��_hOP-�.$�
�}�N2��޴�棣+<h��K�b�]<���~;�1_vfĎC0TXk�@��Z�B)e�JF��j�+3ebBD�� ���,Z?a�p`�����2�>�o;�N��*��r�s/���oc��2��\#tz/�%w�@Wq v.�ઐ���]�yH�zM%�F@KI.g$ָ��l�?<H��)�a^����S7�z�|j
��|�����%/&lQ�	ۇ@�J[}�3��@�=�+E�;C��{h�
hǲ�I�\;���u��T�79��I��t����<ML=#��_U����
���t�uP�X�t6����x[����\PO�%B<�p��y�'J�m��dٙ�f�>�<alH[�⢴�Q!��괤��oC� ��(�����Vl{����q��c���~Y���)���mH�?R���}��]s��d ę�+�(>w�x�����R����e��8��2j�C�3E�;�,,�e+�V0Ϣ�@�#�� �f|s�h�J�T��<�K�bDА��'�5�[_����Ѧ��+e�Z6i����)�xt��;�ȒF!�W�;'�H�B���$bA-ǟD�^�{9�8V�D��Cd(v7�T����}��V�h�e���֕�eۑ�k#4"���T#�2.�#�K��Ջr�^3�%$���׻�8��[�Hݻ�h!ɵ��L�aO!W����;��W�Ai�_u�����|Lq�P�V"�(H��DB�3��l�aзV96�J��K���3�����Bi��"Ѽ���p�Ew��e��<���m�I!�Z������Pp(��33���N�TZ1^�k��䒜s;1���%�����
�`,s�]�⫃�������e�K����W=����Ƅ�VA�+�xZ{�p&�bZ㳃��U ��\�O_]~B�o��*l0T!�}��/2r_�WO��;�!߅�9ːs*[�&%�~�Cg/<�����z���1�Я���i0L��l��ƚޮ�!�ul[?�C�(� O�I �M�Ҿ6q$����+P'��&5�أ��e���g�	�K��ˉ�.�_�����9�9/���P�η�(VW�y��9����y�?puTB&�M��د������
BX7���bZ��'Gkm�E��$�?X;&���2�cI��,�\9lU}c�g�np���m/�,��Z���W�����=�l®:�{��	j{zT3��j��u�@�ݓ�^�*�W�&�jcw,'�X�ֹl~_�K�}�jw�jX)U2'��OJrZB�����Q�Q��S�9���.S�\���ƈ|�/NM�daTޱ���w}����!���F�I�'c����~�;��qKf�V�����;l�m�� �@�Ro�]�qL��%~�k}�G>� m���XZM�3p���`d���b�z:BP `�>��2�y[%=��Nl��4;3���9�1�f���i𱆽�W-h�R'vn���g�ڹ�d�&���-#���@>&�P��T���ט-������R��n��>���w;t�����J�]0�Ng ~U.�\��A��$�x�M����>9U�َ��\����+���l�����E�M
�%}�~?TQmya��`(0k��&�Kn0�5���]z LV|塕`8k�����6�E
���h�FTF��mwu��̠z�WH#�]����w��3_Hi�^0|��h��/5��_p�Z����J�l���@�z�Ur�aβh��\�E��'F��x�.7@�$�������,��j&�зK'�yCw��4]��6V��Xa�P��Г��ܐ ���'�k�S{�����{[�uM�γ�'V����0e�m�ʦj.�^0��w�=_�3`oE�F,wXL�������Q<���.g��L��~O�<T;�l+�wu�	0b�A�
��7C�~��^-�D.W�bLܦ����.�9z�}���i�5ђ�Ue��d�&'�՟/�#����8��J��|�Ωc�Ǐ���a�u���.�q�.�^���d(�{5����f������m��1P�$�z�L��%�j�r8D�K,���L*���$�����u�������xH�`G.��� �|��/� Z��k'��}���m�2�G(��UTIz�@՘�3����4��V�L�c���Qw���U[� ��!5R0�K���y����j�}��{��YԘ1�Q &f�������Ƃl�z��ggtO�
Ռ�NQ���M����>�n��&]��d�*��=��
����Vb�0*Wn�?7����F���&���X4��c[��2���|*�X���s���|�	�����=��{I�ɾ\'�B����Vx�璥���w�)7���.��}�~LE�O�cl���x��x�*�]�ϞA�7[։n�H���d���R�Z�"u2{C�kS*?ǖ|2��t��q�թ�L*z�ǜ.rmŢX_7�Ep�3\�U&�_��;�����hHۚ-������I�o��G=5S8��C�x^!�싏�=��q��B$�!{j�$��)�Ȍ����|�	4O��@@`KZ���b��ٗ!��^ǅ&���W�  s�$��=�ͩ8Z3hhr�L:G�:e+�`�F�����h��X1�J:��"�0ڔZJ6GJqt��x����wwQ2@<�}P=�ԭ�8s�\f��k�cO��B�ߞ���#���w/��ݨ�4�Payq�[L�k��>Y�������%�K@������kKY!�v��C�y���U����S&k��I�0�#IO�!��yL��J.vko���z�*>�F�HkP��J����ݑ��.zc������4C����r��pU�n��;p7��H��� ����s-4���8�TU3�!��j��][N�IY��7��(��LC׸H륧�Ҋ���]��A��L�l��_�>%~J���"��8��L��Z�<�g�1��[e#��2{s_-�փ�x�|�Ev�j����{�0Jr�#��7�1=��3G]j8Wb����S2�.��t!�]0b��wL���7�(-m�	vM��|ڐI����p1����z�6���h�������8Z��On5$�®ڔC,nt|j�eF@1@����C�5KyE�s�=_���2���Z���I�uDS��C��r���������״A ]g��t����H	Iz[�|��Ș����"�����1<$y���5Rw[:[ Ǳ�`�۽�����	��@�h1�	F�a��!�Y�R�6?��7�W!?L�&��/"��G@���dKK��>���w
	CO��+@�Hɴt�t& �O��!W�4���eȁѧj�:��Lt��~N��0)�(�U��M��o?��3����Cs~Pv�����J@We��*NV�{V�/���a;bz�l%�f��a��.]�Њ��#��Sح�M~6�"x��!}���z�49]J����1�r�#�r����0�_�,�2/�S�������$�̤J�ɑ{Z쑇�E9�����;劾�]RU�^"���
Z&w�;?vZ0
}���y����Ĺ�� �˄����2^^�r�N��n#�1ȞR���OM7#|����:�DV�V#�GTo G"��g'��X#,.
��Q��F$��S4a�*b�t��uZ�Ļ��Lvmr1�npb/�>�ʅM��u5�J=&+��g���߃t�݂=�_(��"��m@L
Ĵ�w�*|��Lf���Z\��	@�:=�4ݾ��6���ҏ�Er4���83:so�݇
8^a��(�f��ڜ��a����Z)9p��F��6������Hu���e����J�}ZZ���c���y	���9V	F���Ue���M����6*v�?|�9�1�5Xo���DXnKg�ue��ɦ�x>$GfR��4ɗ�pB�����sA�|� �[�7xae��=��.S\�O`;qʣj�~�\OggU�+`g�Xk-l�n�FDoS���yWXe]:~c���_+c7}u1�ʲ��C&3���9��;����u��J���׏y1����s:@�� �8���X�f(#�T2R�}��Q����?M���yo��p�v����2kz��)�k�Ͼ��h�oQɲ�?.��\�(�I�9�c3`,���$=������){:@�8C��� P�wo��؛u~5�k��Y�l�/;��j�e�O�չ�ܱ��5A�����yX�
V�(�zW�ˇ��[��NЉ�>=���r�> B���_3$����娊=��U~]�;��D҆�B�?Hm��Z�3XPw.�I��/��຾�
zH}ǿ�����N>���8f��Տ�������}��+˺�e�͆h��rZR7&�_��N�u�=h����Ӓ*�Yh���,�f v�	.�7�RR�U�9y�m�^�U���1R\���)\�$%������q�"G+%!�����,r�:paJ��w�����7o'�Z����)uH�i�"$��w���RǺ&)�JVuQi>�����=+�p�t�V+h{C¨� .r�����������kB�3��}#��kE�?���>��&V�F`�܈�J��1�A7g������s��H�.؝�w,ZH�_�
���vl���$�!W}��7'��i��Ͷ�囶ݐW�!�ft�Q���r���W�D�"`�̲�qr��v���5G��Pˎ�E�����b�Eh��b��Ǯo��p��-@D񮭕�b��{B+{���K��o��6EzG��Oن����؇�'���������%���w����C��c�7���8\�*��1�0�@v�	3D�ݳ�A�S�Rej?{8��1ܖ(ɧ�=�D�L5!z+�ۖ����5ܹ2
�������R��HJ��\ r��r�>�+���rEf�'������J_�q ����_Xe��O����D��N�Ջ��E3�N��H�p�|���k~6�'|P��7��Q�}v"���^���.:I*�+�9���M�A7$?F��b�F�ec_���uJ3�@�*�K�BN�V��"�#`H����6�65I�{��C��'����>e��#8g5s��<��4���	1e�ϩKG�<�dj�cv�X�^p��f���":���XX�+6��Vc�\h
�ĥ��������7�^t���$;���us�-�QU�%{uz
`1���ëv�}�$牠f�{��N����.J3���W[C�j�Z@>ki�?C�{�Y]�r������Q��Ì�RX��\#%\�Ф���s��L5�Ց���m�K���0,R*=bl����[�p4@JXx�h$<��wjr��@*"�ϯ�>�4ė�\�< :e&H���:���h�6��������f��u�J���(����+�1�ڤ���H N�B� ��r+C*�r����R�d��@�£��}ʯOlP� ����y�"@�w�oG�ݵ�{����+�1;���ǣ�޾���.�4O`Y`����n�R<Y�i�l>��tG��f�J���G�Z���Z�_�;�-�!�.�&aZ�d�5��KH!X�$��	B1<���QE�B+�H�s�juk_�ɦ���<����q��9�3^+�^N�Z`B+����Q ��Ӽ-�y3`Tï?ܤ����YEF�W�b��aE�?�"���I�dCO��|��zU��8�MC/��۔'[:e<���Jēz}Jjiկ��B�{�-f�
u��,Fp*��&��<B�}��?UM	�m���QL����}�hTf��M�td���!�3!8�-FgG�va_�:�ҏ^�%&˄9��5���
�x2}�q����AD��(;����R��[���~��r/��T���:qj�h#ȉ>q�#2A��G�W�%�Γ��${;�h��9�HkR0o�Y�G`0bi��Ԉ6s���tP�����K!�NB��Y�ߑϒ��$��b�mO�1x3��9≖�2#K~�&�m�U�E�!R���d��եQ����nF�@�b3������S���3��U����F(�.T[.a;u�@���^�(2g�p��B���H+���ΐ��3{S<K�Sru3F���=$��#]Zͨb�ː�I5�g%&���
j�9��&x�;l?�kc��t�J&����{�>�D�^uL���K�-��)���(�W+�V�6��hNR4{���a]��Yjtu�;���c�o�L����%v<��a/]��c��!'��ˣ�Z��Ê��r��	q�����8�Cۿ+t������l$2�5ѹܽ�43'Bba��f�T��g�1Y���"Kd�N�K"�O�l�P�/��
Ì�P����y,�~��pe���9�+z���h�e�ً!�K����$�G��{A���vv`~>~$$2����$<
�bJ.v%��0��y	���E���O�)�ns)�4p`�H��`��sk�+�4�\0�<3�$>�p
I �8T�\UW�rOl��*pj���V�Ζ�;�v��l��6�U4�K�����m��VV�^��WoS���	�L�m��S��o|�.�{��q�e$���={J���'Rɹ�#�V+.Ɗ�ϟjXu���^�%�d�ή��Y�
��~v��&T�'�r(�3��>w}�AN_j���K��.�W~�2���=�3�;|Ȕ�ԦŐ��,gaWߓ��<���O����z�{�[��Inۥ��zs�m4Y���7�<�f!����mt�{Y_x�������<���NI,����4�}��귏48���5�kT-A:d�i�/V�ι�u��E��i���˃x,�@���S;��gk�e�K1u��xS�<˾��`Ǯ��M��@ V�l�7�e��͇\����{��+�
,q
��X�����-lIA@d���B�KR7���]'�9��z6�d#,&A'����K�[2����lQ:}n��hBb����5W���f?^�T�I܎& ì�+3l�(��];u�=������3����ns� �?���N'�_�6hX����9<��G_��u��*�d�|��0"�J��	R?%�8�:�:�E9O�s���L�h�T/��ov��.v�I.�a2��5Y%�-��lZɻ�^��x9׸FtT��1+��C�m�s����ŮU�cq9�1�Pei�И^�u���7H4N��BF���̨�SǰJ�d�/XR�ߤ�9�7!��(��Vl3/ë��A��b>հ���#�>���#��I�~�J΋�^?$.!"���b�s|��1L�a�.g��꼚@�Y�C8�a��*?/�&Y�t���P��$ϟ�OY��v�d?S�� �J�
Ai�"�cY�|㬞G^���<s�L�u-\����.oo�'��'e<�\�P� ��z�gvFg�jG�9�Q�Y�I�:{����ý�r����^y�wM�$�O^�M�S���G.?l1,����٢��x��~'�c3.���іK�����x_��f�+��$X�}U��������O�>I0�T
��k��#�wᎌj��p��C{��.��^��)$1�]�3�Jf��Ւ=�T`��e�P�~s���G��m,��d�|y|�j篍h�=)k��#��5Щ�m �:�f���;�,�����7��M
C��uX
���
��-g�r�1�����u�����!=�|o��<A�kp�4w���cA�S�9���nG��1<.���U��Ղ�tx �
`���NrUb����U�_hЬ��n@�$ι�P6n���E�2���":�`/Ww��Zw�@�g�\a��xɜ�����҆�J�	QP�K�w�tH����J�/���ê����V?-��ԚE6��'�O�~>�y�:��;A.~2��r���Y^=?p���d��4`�����"��9�]y	���9���{_�oO�TLR�L��!a�0ڦ��D-�g��Y߁�C:��z}ϥ����^a	�s�C3�|�j�ۗ��i�b��V/��I�A#���rk�zQB=���|�NۛG2L΃1)�<ع� κ� �6�Ιq_�(�J��T���Q�� �(�߳줣C���6�ԭ+�Uݶeڧ���!CΥ�=��
 k�y������lt��27cj�Fl՘��}�i#���X�W�y�#�������VXi(��c����"Cuw�v�y5h�1
|7>^6%���]�_��07/�*�)�������ߎ�C�@`������ja'}#��]<!Px��ꙝ%�&���@;�Z1�`B�$ ��L�|5��%�X ���J:��I+�ol��LE'ݞ���q���T	J�kjAL�Ŕ6V�a)����I3�~A�wD;(q����?,��mA&`#f��?̱���f���ji�Fn�p153��
r��A{���R4u�X� s8�b7�5�+Y���ԛ�4\�Ύ|ث�������═�?��T��ޕh�!�D�?��S��lM|%������6�O�C��i�,�,�|��xOD���r�d�����-������W���S2����h^�S��"��/P��'%e&�Vo�%8��#,��31��E5�?���=��e�I��d�d5ȱW�������6��������Q�F~:� #��ty��y�h�]�gO�3Lr_�a {���#F���8n�K�c��m�ڐ�'��l{3��v�s��^b��O��q�X�q�>�U�����%ϗ=���5:��#Dܷ��f�I��M�	g�����f�ޱ_LT��c���[��h�T��=��t�}�	-�SS,�@ɂ�M&���$I<�nh˃��i:�ɍ���w��P�b��5A�͓#�JO"�)/L<f�J}�^NU�w�Pv6{҇=\EC~������w�B��4s��j�Y^Y?_GՒF,���������K�$��3u�C���>c4 �E����U�ӟ͹S���U&��+B���`&�(�HO����6�l:ֱ��i8���Gl�0c�)��iR��Kɲd��Q���֪:hf�C����/$�է��,�R�>{�Z��3]�G���˖8���b��������tA���s*����άMT��a���P��NiY��9��<�hR���������g�Q�#��KjaZ3��JP|�f�c�wfH���a�oF�ΦD*�A\ _ڕ^	�G�U�^ٓ�TRޣ�Wzkr��	g<>g��x[��&�t*���[����_z�V�aX����P$��y�b��X��?{�:wD!�̻3S���;u���?$��ej���G_Z�T��>�����낒t���F����Ƅ���U��T�uz	��Uy��n&�9�nu�~���a��Lɽ��qVS�	��ᮯ��tv@�i��?�����EU�����̥�\I�����:��ogd�ʙ'��曖���k�+ü!��	�ܷI1H��v}o��JI���>?w����R���!���A�2#w���&�|W�O]���B1�vc�`�9�K@�߰:������q�vJ����8��p·B�9��48�ォ�\΂�/q����k\Ѣ`E)���1M��j�Q"9y@��WM�u�ܔ7Č�zb��u��&���>����l] � NE�N���
"t�d�Na����AXSSjSm�>�3��[�Q�M����ZO�$���`UY��Dw7^ShQd�8�D?��h��	��Rla�J8#g�@��20��>���p�D0�[�x�D:8E/�%��HBP iIL��3^�_�U�3��>��ߨS��`BYo�\T`J՗�� sv?���( ���p�Z����L�i����6������o/��ͪ����n��t�ʁr�J?ɪ��=o�h��6Ōz�v�+�4v�����؞�����F�:��1 ��P<���Ew��d+�y��E�����*��U�h�s��hN���:�=]��ݿ	`���O� "�w���I�R�����_���_X�������m�~���"�=�N�88�-x1�B$� l�r�
���`0�ZiM�/hB� �)�-xt���bdTj�$���%���(���aG�g�Y9���T�>��5�f��ZO[��S����'��|W/�|�ٞ#��.b�k�$�íU����_Q����3�H��������e�=�C/AZ��+9h���p1G���ܣ��ٴ����WSӠr���y@�E�����
B��,�E��{#��*�_C��(�6+�x]�~SXX?�.�R4��Ӌ��B�͆�n��;k��WC�������s�B4:��R벝�*Zt�i9�,��!�(;��v���4��������u��b\��J�F2�2�CȇhA+7�@�R�]���q��a�N��� ��=����<�%a��d��sݬ�S���V0�	����~tX�^��\�T���o�f��P7����~WA�D��ַ�b���jo[�ui�}O�{R���3�����I?��᤮�'iAà���hS�rU�=��	�+ۜ����ښqR���I�0pG����Up(�P�]�W��0���N�2��J:D' 	��P���3�ߡ�ʧ���ö�X���Qj�L`��9Q\������%㪼`s̴�����3lW�Z@e����*PaBy�*�[���Ba���/���H1���x��o�bN�����];[�ʨ�����9�ܙ�'�H�ǳG!TES�l�},U�3�*��3/�ñ�?�����מ�U/�V#]�!4F��>��c`0�=�2�,���<��a�)�h7M��+*����q�碊V�4X�����3$�V�b��1�-��ý�-�DV�K�ZN'�}6��$=�ӥEx�qt�]& Yd
��c�0bZ� {�!�A���(��J�,�/�kTx�z�\&ݑ֋�"��.�/��p	��k:�,s�X�v(���\r2��&ZK�`9FuݡY)������ ��Bzo�˪�4��ٴ���[qJ�*,~��8#m��a`L(K�-^Q@���ծ �rI!#�M�S�{���E�S
/�L�5ғ���Ɉ��_ �&9*^U��t�`�����k��}��*�=m���eҽ���hk߬$��K�����Rܟ��4�J�h�Fl"I�s��UW��o����4�U��^J�A�R�(h7�0r�(��(t4LD*C���)f�+��\+Y	}i�� ����;�1���/h���U��0�����p�C,�G��R��9��&,ga&I'�k�%��|������P�l��>>M
�i�`���i暳wd&/�`\Mewy|'H����R%���{�G�2�<Y�ؾ����{{G�L~?ƛ�*�e���|��f�����8o��8i���ū�e*���a�m��ر~ʻl�e�Ir�ۄW$̼a>����o����ь�	  )2t�%�DBݫ"\n����;��+i��,2,-��<#؛D�O�UK)g��R���끺�iެT�˱�����b鋉)O���>��8�eX�$���Z��s���H���Q�:K�}��}�!�5f���pn��>�����n���Ŏ�������}��s����|@���N�����#9��=�l�������o}���s&�5���6y���z���4��!y<�T���	�	L-P�}�T8#Jz�֒��(D��ĺ@G!a�p�VO,0S�ԏ��&k�}W~a�rZ/x���i��A;�y�ꄒ���r9�eCn6�'�xs9�#�����	&F���Ti
�r���X����@�^B�Q0��G�Rӹ��b�F��+h��Vm��U�	�=�	�[f��N{�x]X�c�̭e�^c�T�Q@E����ܰ"@
���܉�R�%&z�z	Yѳ��d��'�6$s��į����9���H��|hE�b�gC�_C�h�c+M	��
����� �!Ş2�#k��d�.�v��K6�$R��,Z4d��'�z([)S3 �����FO��cqzV�����P]Hۃ��r��o�H. �a�Z5{�]B�"��ɆXxj��x2��� t!;		�x����̨6�tw9��ǈ��Q���6���$��n*5F6��.Y��O��F����mBnT�P�;c~~����
�+
�K�1�ɫf�UiK��!�|_��F��u�"#TǍ�}Nb]�Iψ@�a�R���͖�|�j^�9�l�f����2�K!��/�"<<�.S�����G-�z��HX�-d?v��Z�������߀�N���|ی��q�VL����[(r�i��E��vU�qr�߃�
e�zC�9�gb�o7�����+��KZDqaW�q�`n�E)8�(� #
3�P�cU��CۙP���a%��{�^��37���S�!��6L>���1�n�葌C�=Hji��A�?��9��	T�g%7�K9�r��Z����Ue'&�s#��yF^�:
L:�^��j��nvM�շ��4��k�í��j���¼�n(��+�'������.
�G�칩(��f}Ά&�;/7x����[�����Ļ��Q�'���	C�<5/-�'��ID;�4_T�X���R�ym�\8@B���x�^��*�i�l��n��g�o�Ŋ�a>����K���M�=q�ӒW��J,7(��]��4N&�{��~_�P:��s��V���р[���1nio˘��rq-�땮������K)�p_���t�+B��n�&l�1\؟OF��Qʊ��Nh�[��I�r�	�����t���^�Ӷ 6S ��I�;��gOD��2+�Xc����T	N'AM�N^��e�[:��1�1�6������/�Z��%�����,>\t��]��@!�3$�Z�3(�0O=s���S�d�:�^L���,�����4ۂ���n��a1�4f�R�� Hq��5����yJx��L��i�||����rS����t��̪� Ӕ��d��BۧhsЅX������͈��ӱ��=?-��d&�^u��9v�Rd޲3���[| ���3�1��Y��d��R2���=��Tt��&��̡��7�vU�7�FMw�z�` \�e���Ls���T�R{|��{�E6	r�E��Pź��D�~�'���R�}�F�<���b1�����DAQ�DO)�p����%�> _H^���)�	��h� ���$�b�,oMA{U�D��wЭ����nV�O	���a�����s�5;�`COL�91�����Ч蜃X4��Bk��ѝ�>�{������\G���0�x���&f-�p��;��Tl���c(�#$,��{�n�e�R}��l�;7�k��7���y���U��[�?��"�%�$L�h�I���fb9)X4i�\].��͡��/w���������s%B1�ǣ��q:c��q����v�����N*\Q���.����9y�V�B���&"9����	k�j�&E�au�1���zOKcvf����䱡�Nit�6�
�� ���Q���ƷG�u������"#�R�D���a;�)TM	+��kv:ȥ�`�Sr�[��pI�o�3֬1�<���Ch9E������g pU������U(��jD����R���&l|[O��T7���}�r��D�j%�v�o͌�H�+>/�����]�q��b�l��8x8�ƃΌ�?2�{K]�<��rɝ���'����G9�)a?�������Ȝ�����s:ys��goS��Y���,[�I��U���A����Q��s�0��h��)C�9����3�cQ���v� ���;��L���X��W+.n�\4�^���H��N,v�,y�0b�g[�o��E�}�,;�L��5��#*��`��*A�q���/���r���C��a��c��ٻ%��z�+�U��{@�+��C�N��pal]	��ѺgQ�\_���qq��J�qrB��8z�$�R�i�l�� (gf��a��!��^P����$5���w"���(���	��ɉd�6�|�H�|ok���g�U����5.�h IC51��O�m>s5Å�j��1�n����;7�Q�5m�q�)j���Wk':0$ZI���D��ګ
y|~��lU�+��E$�>,�.Dm�h�Zf��Z�I��J�x4�8����;Ĺ�'��5f�b4zs��������B�I��7��~�*��:l��v�P}���$Z��k(�b�ơ���?[m�fCb<��+�����bǡ1:i󳫲y�"��yи�8U�\x^bL��n(��0�g�px����)�T-s���NR���B����?4{˦l���9�<~:�Ɂ[����������Μ,��q 25�#Ua�D}�&�)�Y/�`n< �Є3#H��?nIi~�,�0�Cx�;�z�N{u ��`�y�%�"�2AW㴲�I\)%H�g{/틼�}��tƱ�[E:؂�bp���崗���)�tt��G�cҦ��6I�~����4�������w�Z7R�K9+��&ESc�?�D�68�.�2}s��@�t���}�m(�@���*WU���2�UiwqN��B�օ��kX�?����)�Y�K��uR�?3U�粬i��ck�w���y���O�.�S���':��e��B
i­�J�~p�V��Y�)a`ٲ@��ǻ���aNX�^�<�/
۽,����-�MX�K��)� ��Z	�	��Y�&�לs��$�� ��^�_Y^���w��	�5��Mu����^��홖~����]Z����Qk��{���~��H�aP����"��,TTt]�"�ntP�x��)+����,J��@���A; �����S�8|�p��A����֋hH>�9����sJ7���-�NO�H\%<Q��N�)M]��{o��DBf\tu��.jyY�b^���4/����d'��ʍ�����I��N�������p����t�~��3�Q�Huz`�9)�s���?��D���֫��n+ɟoW��}�K��8�Ma�ֿ{�[�!���p9�� �"Q\���a�]u� ��r�PJ�~[�f�R�w,�X���/��(]{��Οw5c�����ЅFT�Z�gL��0��ssЊU��)�O�^5-a���|u�QC>�/ş�g���J{�(��:��Dm-����#/�t�=�X�<$�sA��ȋ�Е��V�Z�CG���*����uym;T�J�耉ػ������re�7�Ν���o�� ،le���'͡Wp�Dc�.�E{�-tݮe���.w�y�J$o6�:di"���8m���y�}�=/ౄjm��y����� ~��U�,�5�iI�.���O�r'6 0I���k#���ux|J�����_Ú�3IDS�RQѯ���wm���lŉk��Ku�\-[�g,g��F�Dtq�@���==��}�Ѯ���6�%�2����҉��}�T�֦%"R��W;[ۭ/�&e']=�@�0�n[p�ů&3ҙ���,x:Gy6N#ۋA=]�Bz���hf��b3�Z�0���1��2p� 㯝�Y�������������`�#��$��5�7�����z�y�pMrz���k�)���P���Nr�>g �@{�V8TY,�8�#�i�4�ʹ�J�D��rC}�y�$��x)�o)��\�O����V��#�)iҵB��/�#	,���}T@Q�;~�q�h�F�5�rO��|���<�I� �t��|�����g�����y��ۀ �������I%r��̖���T]�F=
�t)��,��>�Hl$�O�W*)�$K� ��;��W|�<.o �A��T�n��(NB���� �)��E�^uN�Rm%k^!A�v�
��3j(YQ)e������M��0M���rk��ՅnC�S�׃@�B�ED�BS�ᡱ�#�3�Rg�����J)�\��@)JY�G\��؉y��_ۊF�bحY�0TwnЏc.��G���~҄߄	 !򙎬k�3�[�M�,\���X�Җ��v���o��L��Ťo��_�_ݍ���p�(n��m�(�Ǘ�>��R�wM$�QW��n�M�#ieaH��'^����Lg�d�7k�����'^z�K���9<??-�m�H!�C���*
r����}4�n�xCn6m����f0�%bK��O��X&�n�#�}�l2�u����®��lp���r��,�h��5/��F�Ӥ�3_�]�wlnwS	_��ªE��K?v��9J!�C0�DJ#f�
-��s�^�B�d�3�W���ד5�{+��8(.f��7�����D����1u$��e�>�,:�X,x��*J|�L��R��� �v�Ǆ�70%�S���`�&�J�H~.��yS@���PnsEX�PRmn1�	T���^�L�,<͇�,oҽ�߽ֈ�A�\>%�<���M����:Ia>h�8?����2}p`mq���ȯ����S!�'�{K�Y3l!�|�~�lˀW)��¿�(�'��9���z�;�cԕ!K[l��z��3-�G�aD�'��ֿXZJ����1�ʕq=�H��!�"�1J��w&]�s������Fw�DM���н�e�`��JENs�{���u�*��S������=�F����{�AZ�WM�=?SVͣY��\GZ��j�;�� ��L*S?��3�`�$�Vn�G�h���~P�Ջ8i�����&�`�#x��3��Ib'M�K)��� �ĩ%<V��.t�O��Ecl� &�ܗ�s���3{_σ���>����Ng;j�;�� �p��B���~���?���;�����o��FK����i�t���a)-��vs
}����$~ov�U�~u�cY�a9�,,|3F<��7`;��b��7ߛ�t{��>́Zl�H�<t�;�+leʓH�d�8g�5|�`�9�\V��?E�.[s��&@���X�O*�:9\G��·ܪ�
7z2���z)�gz�ø^�l�������6���q�$/SiIf(?������
�K�%C��ǘp4IpNZ�Kl9G������Ȼ\s���������[8������/�/���MCl���Bc-�Rbt�_�T׳&�l<���U��vb!��XVj���w�{N짋��O=9��MJ! �0�kli<����B6�]�9�˹�wG�/�:�E8�Gg문%vF��U�,e�MKp�Gԁ0C�[%��C�����H��D
�����9���V)}:�� ��l9mx�Ʉ.�.ё�U�MH��3��,bB_ �w|8��v�#a����
D�uT���P	��ˮl
���@��~'_ }g#r�=�{��[�G�v#���7KV�-�~J�2Ǘ��>>)p�/��C�DQ-�?��?��!Bc��p��1J=����b���EAAe�ӱ��&�Df�PkE�����ug�Q��K��+щ%��$��Qaz�;DM,�X7P~��.�}�	��cg�l�)6a��+Hv���X�^i(g�'RL��$��d3P�_ӽE�4pU�,7�pAE��~9�`<���N��Ve�H����2 ��?w�\�Ǘ��N��CF�&��?�S_3?�q-��aT]��.H��TB�����<��ҳL<�HLa~�p!��7����Ib,*{�`�9���H$[e��~ɗ��������V0��Z�Ö�އ���h��j��*���w�+�O�J�k���dy�ŝ���d�X�Ww�o����ʠ)�ྼ2��a,@r�����<�qu�v+�V����&6�����ٯ/}���C�3~�4�:7	0Z�����$����4m0�v�~�g~��rm �bf'�E�q|C�������'�'���$��8m��N�i���0M��,gM�fE-8�u$�����0�݊��*�A"�i��԰���*��{����VwM-�/�ʜk��L�|�%S��h~��3F��K:�JX<����­�q�)��5t�3$$�f��g��j̣�V����2Xʵ6��5vf����9t�E�Ca���x����c��m�qaG�j{����lZo�m�!À!����h{���5��|5N�����g2�\}<c`=��/�k����9ώ}, ՚��UՌ�N�暽��髙��X�Q�s8I�}c��9#�r�p���0^�[}�5�m|�$�9�9�q�/��]�F-����M>��A*]�g&��r�;2�ඵ���C;���&Z�n�@ީ���j�u�1�nal�հ�O7�ӽt����j3B;#�����:�UJ�~���S0Cj��LG}_��|�P���Hk�����l_�v��ı�]}���p@��2�kp�Ocu����5�h#�oꞩ�ڻpOT���lUK4�1���HF7����<��2k�*&<�Ru���{
�Z���X�����R�C(|op&�������v���~��f�X�?o�_����\��&Ÿ(�g�}��� I+�<e�o$_é$���M����%�`_��Í�kG�FT�wZ�N6�SZ��ϐ4ѻ�==[p:�Ч#bD&B�X�X�TJ�_u��H��*��*\�0�J[&�B�e��E�P8�ǀ���N�+��k��p�x��Ґ��dMx80��)�;U1�G���"Y�޳�����N��N&wP��y<BWz,$�n��WL�kNU�/��{*s,HFM�ep6��{Q�aa�ٷ!I:�V���`�����Z��X�6�D0�gz��'UY�~Q����YO��|�+�,"�"w�SF��ѩHy��  :�'7��@?����d���{�E�G�# ʬ~�SO�Oy ��՞�MM����ߨMgv�t2<�CNt0Z[e��Ji��7dEI�Alt�й�z�{���ϫk��Ы+zw�b�Ӛ�wrU�~����y~��nu?ywF�<J��M,��i�c�h�k�4-�:�&8�5*l^6����4� c%����s����J�=�jdE��V�f�|��x�n8�7�G#�Z���rK��ȡK�fi���(�
;[���9�օ���
����/�@�ct��
i-�f�φ-��|�0MuUɓ��X�.z1ΰGDd�d�q(2�欜^i��xU˒ɜ����=����t}g���v�K-t�� S"p�E���9�i�	�?q<��������!�N�f�0fh������L�$��w	$T�G����!�W��^%�|����A�hZ�-P������i"�03���ħX�������5#�9�
�F�dE}�r� �!8��?Ŀb�-�3�d�������?֋Oͩp��y��?E,�����Ь���=jP���W�$2+:	(����\%ODs)>�8���]=��ɣ���YA	��=�9uH)�f�ϾL�݃9��@�`���3�WAom������2���F������t�c6��I�(��l�u�����=�ꪑ��3A�ƕZ�=n}�Q�dE���{4>�+~�|���a��?��_��뺌��`���	��ю7��3#���K�&fN����ّ����d~{��
�f_���
+f��|?e��@z�s�m���K��f�EP��M�e ��
��_^�[��S�.7_�Tj %��w�M��:79�vquw�X������h_��l�]�Ԣ�r
��� �t��QJ(+(��K[�'Z��-!C�x����"���%���2���yՊ�
�m���Y�((Qb64G#K���O����>�7�� ���YY���bê�ǯFw	�]���S�J����-t��=!�&8���b������Dk�{��r]K�nu�ЁL:�I�a���|���d��b6M�b,�	����컏E������=��n��N֜����a��͋mާ*=�R5��8~�����`#?�K +=�,'��0~�C�̏���Lf�����H�#�~��S���2��{�ɤ�t��{�-��獸��)�/�*�V����׬ ۬��Y(�J��4�F�!�&��SRi�#���^��8�Щ�Ɔ$��ax3�u�2[�F�|E���Q�N��g�U��։�oW�I:q��Uy��|�n��z��dt|\����zT"�� ���O �	��ɼo��X~�d2=��B#�y�r�nA���U�����
P�jBZ�0��i6Ņ�R~>�B�k���O��;wV��Eŗ�'���^��P�q�wH���+��m�	�I�?F�Ji�E���d��/���{���H�8�T�1����a"���ȟ�aH�9z�祹���v0s�WOČ� ���\�f�����#���Ǔʥ3��$�'k��e�AOܺJ��0�h%��	���T�y���L�3&˩���,����Y��֥��[�4�S�����л�Q�5 ����`�Mn"�b�1���?�Y��ht8��g��P�����G0��x1�a4L��a��ʥ9ħ�`�	V���k<�`�Cz.q���D�U�˼���] �����@R�[ɾ���y�����0���d��kSSڣ��%���P!��|y���+�@"��۹�^B2��\#`�p�\֮�iww�Vի���?Q�(F�����S?��B�	%���;9��n��������A�,N}���W����{���s&�e���c���1(3��Fa�ߜ�N�~a�P�O��Gdpgq����d>K.�Ѱ��"���-1�@|��D���Z��k�9�ɣ��B��F/�b��6��=�t �R�dWDC{/��?��]:rbX�?+��s2'(< �����������S6���?��0�W�i-���:��%�~y�A�R+�&��4;é�!{@�V�sV�A��^JY�|�4�:ZtZ�n�]�M L�~���� �\l6�X��𜛠� �T�K|���3����;�靔[���֮�j�q �1D��zf�p��\��H�S��j��s�Xf�ɍ�_.�o���0$L��$W.6}�"K�zL�"���%���t#WZ��faWd) "�E�'$���2��#.�7C�`<������Ѵ~�W��R>\8��u+3�5Tw)B_��H4Jm���'nkN4��|*HA2���a�,2u
�iG�6&;{8S	a�J)��G�:��eX�+���JH+3���6Ji�޶���B&�t��B�T�<J,���Zy�su�)�+ZZ�}=����J����簵#@��X��P�x5|I~��ƓА b!�O������i�>�����3Q���'�s�O�d@ �#(���	�?�:��}9 �CNl}�����P��7Uy!���%�ƾ�ʰ�� �k��^�rP_g��W���Ħ[_D}�y�#*�X`�-����}�6�Y2N�&��jlh�:P|�+p��U�k���mqHX�0D��cc��u�W(�G� �Ř�c����4y(	՛"��/��R��v �Ә��%��q�w�� �[h�
�M�֬.��4P���Bvh���i_�?u2&����+���?;���j�U�;�:��vI"|p{l��;F��褲�|�?�t$����(Z�E:��trDQ���z� *��&T�.�X��x[���qZ�	��q'ߍ�ҠэH�^e���ۋ�y�p�ܕm�>e��>Tq�y�_���{��dN�x(#Ñ;aK�Oٷ�p���f�@e_��+V&,^�"��_.�Ϡ�\�͓0as�,�-7���`��,e�f��0�>Wo�H*��Dd)N��0�����,z�2��Qx�H�fh�}V7(F�?a)�~�%w�Qco!z���Ck��B�Dk�*�oѺ�<�!D�g$�vgcL2j��o�7��O����$�ZS��r]ƞ��8�w	�\K/�<ܻ�~��Cˁ{�� 嘅Vc��o~��7p�M��� G�aԣ
h?+;�K��q��g:?\��Ĥ�3�F#k�G�.�� ��C�yi�R��rf�!�j*�.�k� ���t���،��{2ۼ_��(������9 �G;�� |QoC]f��o0��
�~�v�Wk�f�M\C��j �M*�|	����O�@?[�����	���Z����8~�E@a�4���(E2§]F�'���l�ξ���m}���M�W&Pz9�M(2�K	6�ᬆ�к�,���Ҿ�8�J��7V����U�:�&o�\$i ��	ʥI���c�]pK�r&��x �"�����{Î����4O+�����E)��:����n�p_l7Ԃ�e3�'��kVxe���඗�~��*M��y������+G�I���8xX,�����m��S ����p���a2A�jt�����l���I�ϙ��\�~*��&_0x�x���9M�$`u��	��GN��D��X��E`�6�ı��o9����)��D�a��A��l�����^��g�8Pѱjq~��c���h�A������&o�B��=��ڧvpB;7䄹��6T	:P�\FK�\b��[Uq������<2�k������e�G�}vރ�4�Ӕ�X�]mǵM��~I�hN�[trsu���;|���y�Yy�6�D�1ga<+�|����d�z�J�Ȼ�~�2���u�A,wJL�4� �pfq�߼/�0T�0ǈ"￱b)3A�B�]��lzݴ�Dc���vcFޞ��\�Ü�y���JTL��j@����2��"e|�F��1��s�����pR���A��Ă����p)���%�k���#��qG`6�����@s��?d.�,h�&)>�����6�4;$��Ф .v��p�6�Hm�,
Q�� YhY��5��*��O����.�L��%����㪸8D*_[�a� $Y�2�p3MV��wB�>��� ���,9�f��NػL��r?K1��*�ެ[�Y�,��Q�(�Om��Ϧ�ѫI(����W]�J����r�����";���;��&�PF���^ɡ׷~p�?NB�2��K��U��2-�FlpG��?��,�c�D���\$�@NB�b"϶z�ɣ���*C~��~���	;�!���]y&��}u�~�����]5@ɰL&-�-V�0�}G"��^�[�\��jD��C�S�(�(�#�c]���r0�z�+������G��x�E#)
���.����
Kc��Ǚ��g�t����l̔�h�`X��Kgi_Z��N��_HQ�����X�#�=Ș%�c��0�$�PuOX�t�&\�dPc��Zl~2��0BM�)�5��5���t�W\$�/���.��� ^�'͎���j�;v�c�P8�ǀ�sD�') �LG�|�d4x6<���:����[g/KU0�Ũ9�#��b�OBE���;��FJ�l�U�$"�����k[�v}����`�J����ϰ��Z��i�Y��n*��8*�\�Ʋ���$ޣ����HJ$��j*wf�"�3�z��%���j�l��cۂ2�LqRʦ4���
�%'�d��>|*ᜂ?�f�w��б*7��l-S,�	��ҹBD�d�!��
��5X�ħ͗��Z��=���ǪD�?H˙O���eƗ"��CQ����t�@ΆoD��CP*`����o-%�B_�F"�R`�$�o/��-?(DL�ww��t @c�&�0�����d���ʣ.TѤ2��=�aw�j��㧤�d{��7ӳ�3bt��^ *����lR����g�ɱ沍�*S3�� �@&�;���g��E�~��^}�q�,��	�,��?R|	l�7N��@�y�- X-�l י��ݟQ'��������(f ��,Ʉ5S�L&'��n��fAIɍ���#�~���3��H�5�A��ix�D���Z<-��n��ă��,��2@���:_��d��NE (���bOL߽������v�(�y����mz���rZ�PG��k\b`.@t�4{;�-ҽ�?�1�����S��驸<�C9��`a�mgV_��Lo0�3����*c�s6t��9\��������
.K}���oW�{\Kt����d��`f��8�N��S`/3��?��ި���i����S���4��;%���YJn������0���$�����_Ⲫ��M����g��1\�	9�V:��&J��bU�+/*|Y��_�C�=�6�5��ɱ��N�pG��R����$�V��oB��R���Bv�n	b��F��Y	��+�VQaM0"�����;C����j��3f�Fj,��e>�˚��fG^��x7���g�`�9%YiF<0d�:�����O&�<�{�3Pd��pgx+��@WM&Pq9���-�O� �]����%p�b��}��$B�~�
G  v�0��y���G�}��l�r�/��.,�EB<�z@tQ�}��of/6��7�?
�����;�%W��l*Ä�3��?N�O���)z댸{���Mإ�5Z���k�����Z��ܷ8���<�	Α�@Ƽ��̟��(Uk��k���uo;�
�l=7��(l�l-��8T�!+Z[���^p��N�K�:˹]'���F��2zv�s�V��{]$�Jɦ踾#k
�7nɩ��!v� ���	u�q�k�Bݒ��X�K��$kٓ�HL0��~�9T<i���A�A�`d�?�_V88�#��9�]w��N�W��h-_����K/�x'�j��j��߼�Z���s���Y6�� -;����^8Q�X�DF��o]�*��wU�+�%�����Ld`��p��k�]L�N��%��5���f�e�u�iq7��t���k\Vۋۦ��z~)�$���g�;U�|�yR�I��쯉�H�G����m$@���0B%FH����Ȑ����]�M<9^e�r�1�B53l�w��
u����%�@����=n��X��뽜22)��at����#{�C�����s�c0�vuj�ّ�C��Q�b0������?̲!���lg����LH;�-�&�����J ����^p��	��O��%S�8�9����A\ʪT�#4WilD����_v�QӜg��������	SO,���$�����$[���R���փ��������w��
��h�F(�No��9��8���.,�-�Z���+����#Ƹ?�K�U��RK!�?S`h�2��c��T�3�q@�a�����`U�ݣ<`� �Y촊tԈ&Jw�fx�JK�_�O����4y�Yj���^�k��{L��6q+����̦>�_�=h�[��b�^�́�q�{&#��Bz_�dv�x�G�% u�ȎY�W��@��e?��Yk��Se��V��S\ʕ�8K�'8������7�G.��eXp��OC�<���B�����3������@�ߡG�8EF}��W_�Ʃ�@b�o�9H.�!���Ե��?�V�QR�)�8ĝun��9_��@.b3��r ��������o�E��ԅ�g��L�vo��&<��9M�Q/��z�����fT�:d��l{��G�1���d)19~hҞ���e�mVc�C�}���J��������I%�p��F��n��-WV"����3!�T+��!��'���R1�*R�mO���LpsE�(P�S�ƌ�t}E�ԫ�">
��l��wCLˁ��GYG��0���p�X؂�aX�xK�S�A5�H�5����Q݋9b4�q���a�����k���0V0z0���C�<�GX�xw�<@�;�=Â���wyX�‰��TX@��4��_�b�3��Ǭ��#M#:	y����a@ܓ�m>�E�S,��V7���mp�w��72�� �T"�߈�}�U˰!�Tki֎&�gG���1K�h�Q
(�c�̙o
B��1¹j&d���B�I�鿑�i�3����t��l
���:L��V����$�ڙ}������΅j�[��l����_��|��_p
����ݼ�_n4�ݤ�+g *2����� E��0��PchPAי����z��j]��L��R@�2I7.�0�&��kf�B����M͸ml��ՎTbA�%�d���\C���|�3���.Q6�7D[QH��l��]�hX��̹�\n9%1٩L�x�Oc���� ZĨ��]W/F��qLI�Ą֗s�Z]�K���q�ݢe,�1������ld�������;�������퐃Ӈ���L�OYj?�-�Oh��_0ܱrֱ�΅�75��mD5m���3{a�!�`:�Fa��=tT������L�ٞ��xS�Srr� ���F������.f_}�8 FJ릆
|�n���0]�����>�Ov���!�{����Z�W;���N�,ߋ:x��N�����&S������T�)���l�unj{�Ǻ @T�|s��7� Dc뷴6�f�����~-�C��O��^h&3_�h:	�%N�v�dq�Mkn���-�YU�G��C��g�}Q,J,U�f���#/��FI]���)���D��^p2�lk�ʲEꕅ¢��2@Rg�{��P�`C|X�uV���ު_�0&�%��Ф[!���Ϫ:�9���jĩ$0\�r{��)%��לRV�6��c
2�y�h���Du&�6�%1e�����d�:m���؆��f���,%�>pL�l$S�ӈ^,�S�:+B��#mkIi�{gfw����m�hV�[�l�dB�s�	��sR�_�J13'N�=���n���1�<aڍ�ۑ0�p��5Xy��B�+�͕(N�1Ao���j�T���ۣ��fTɦJ�շfe��"�權�[�-q��n(�x�*��ٓ�X^���3��1�g�(>Bxd:�e�f�hQ�������'`���+�Gό��&�-������xm� u�8��=�5WMy�L�1+;w�lN�&(�1���x��S�.���P��~#k��N/������(����4������$[�hV�u�"p,�L�a$��8>O��(r=v�k��Oϓ5j��>�Y�]��
�ɝ0�u�m�Y��Dՠ?Xvp:��~�M�o0���ƱNC,���f����V�\H�`�z^���u�G_zy�Jk�F��F�Ur��F2�Q����q��=ρ"�b�t��Io�T�%�x��|�<~[�'�kB��G�(�>1�����h\t�*J�A:2$�;n�:Yw�K���í�����-�RBwp����:R<\1O�Yӕ5�:�ހ��`,�ы�)�?2�8��;$��)O�f.6��)�yZ`��]P)!
m��Ez7�<T�б�$�]��e�-r87t�Q/�.�!a�~��b�vBtm��gA�FyFq�~x�>�
P�dX���eؤ����K�����c���!���L4@
d���9{!���藋Et\��t�=�M��"Or������� ?P�u��8�I\Q�1<�d?iϕ_k??|���.�95�,ɵ@]1���w0�[��t3<EeB��':]ҖJ��脙$�Q.��:'��=z{�Vʞ(�6I?���j����Y4�L3�֟�<�*�"`��8��f\�i��ʾa%�r�`�{��������2�ޗ2%[S۔0.�;%rV�2�}�C��x��L�����9=� ���n�"sl=Q�/S1���	�[2�FtE������w�z�|�Q���[O�0oyV���* �w#���/�b�'5 �������P	�/��ܦd �'Цt�%���h�{&�q�m�WuYqb\*�|HG[u�~+��B�8�'�A�����؃u�Yr� <Lzw`���J�����%/)H�Y�M� �2�e�lދ����-�og�Ki"��]�Ci���n����r"��a�&)���yL��������S%s��%�U��²��	f��
A
wO-��.��>�Ϥ׳���Ma@���#�� k�o�7l���ޔ�O|:�'zVX�����j+z0W��m�֍4�9j�������㺳k�j漙 }�f�sC�*l�yw��f�Szl�@����߀[�%�M'���al�+.d��> k)|$'����g?ѭiZ1���/k�$�f"(�b%��!�" 2e������(+�~9�נ��c��ޚ.YUq5�-F}ʌ�Y�D�wX('GA�!r��6������/�2S�o��~>QF��|Fr$v]J�F82��$���`�G4+ 7Ym���'[|h��>S �J?F�`4
��)Z�H�h�
>�D4sbO�,vխ����������m%e�`g��H���� ��=��Z�f���F1��\P�ާ�`3��>A�ɪR�,7tGp'�&U�|r�#�H4T�2�de��ݗ������i>qD���G�>��ڿ ����M����Y�Ay�'��'�4�^�pF���G�m�����v����_�� �CI֖M�-�r���r�����t0��цߌ7#��,�N3TC��jv���CJ�̕n	�J���*j���JN�

$�F�{��!x��"ʼє�xH`CE�����Y^��[�;���W��&ekTᖜh��\�6b������2A����CXƣ�m/��ư4;��$tJ�7u?md�}��q	���E�Lj���F�aw^(��۹�d��Å@|����<�i����y�ҹ�p�R\���YG��	����Ip���Ġx¬�$Ó>\%�� ]�YǔL�0]:9����9Ӥ3���w������3�!�P��\Ƙ�5�A������P�����b�}En��:�~��t@:V �^y�Hq�0�+h�~3U���b�8*ql<,=���EӞX^�/0?|�b*}	���J6c"���E����2��h���^9����薨�g�y�/�&'����]��}cx,���y���/KA����A�gQ��BHJ��a�K��G�2*���ݽ�J`�����f��Yݔ������J�S2��Sh�=ZD� �a�?:��{��d=�#@5�b!��qb�5�������wW�2mL�qG�>��)���'�{���!D�:�/��#��gauﵛ"�ݞi�$T���a.[�|M��ڌ^I=�-:	aĞ'�0^�_VE�En���~>��a�8lQ+5����c:��M�����ꖰ�<�����65����/�w4_�u/K��#[Q��<�;����\a,':�m=)�ރ�%�X�uX��-��id���^w��R�g�C���-Z3�����]4��]��7����o������"]JM �gʷ����Z	�G�.��-������c�r�3$V�����Bq.8_)�H�2���z��x�Gh���Ҏ0e��j�iu>G��"��b�6�)��G�#of֙oV(F�[u��:ow}k�#�� �#;��$#Ӗ}�hn�֫g��7ix܌̠p�U���يW�ͺ~��AgE��9E��a�ʥ�Lp���/�eB��3�5�n\KsR��0U�쬁���	ײ6ޫ�0���DTӹ��ױɦ�7}&�K;���F:��`�ɫ�~��}
*��X�;S��-��Tf*ӄ�a8D��@�%�t.};����kZ�U���*��Ԓ��Hr�^^|T*}�sc7'>��\�lX���EH��K�>���"��]�7}@�q��c���*03F@ٌZU�ovTR%��MrJ/��O��m)�n(��W�|�bL���u�F>�cHcf�>�@|ӛ�f��b��y`����	P9ɂ���~
d~�
p��i�ͼ:G�K��㇝��QTOqaibhN������������8�r6l�ǗsQL.�>ot�`x��uf��蚇�@@�V�桝?Ι�/�j�֧��j���s�Ɔ~����;�+�(U��@͍��ytI� ��Ly�fJ�X�=rЂp�d;�VU(W�'X%���S7�x�{id�k#}9T��l�)���>�/���Tt��
.�z弐�}3	�J�	'.g�m|�mh�����l0�M�e=�V�����|3�	���h1��3=�T}{�q�YD��/ڸ`>yi|���uӿ���&	f$��@�@&*쀿��*������}��F��l�ۂFg?P�A��Ã��v�g�	�f���!��ȭ��su0�n {,;�c]�6IKX�h-I3�ş7f1�#E���s,F��1�Lz ���;�Z����tA���@���5^9�k��`�SU��Z�ߟ+ 8���ۚ���B���t]p�݀�C��q�$�dO�Q�=)�2b��������(�f�-�,<��^
�g�Z�F���^�����.*Ϝ 
��A���������[�Ga��p�AHDr�{&gz[��:���t:d>\�J@LVa��x�;�u�!U�c@��	H7jdܾڹޠ��wN�?w�ŬZ�,�h6��ö( v&��|s�ضb��N�;w4[[l p�52��:� 7��b��]���S3b��0��,N@+����(<%�L�蚑 e��I�]���Pr���6W�*��e{<�Ҝ�n��>�ssLQ�@����t4�����=�+�@g*�g\l���I��8Yl�Kb�m��t�H�X��vs�v�Y����-#���+���#�̪�W}�J�2ED����p�0�2X6�������Ե�3��"�2u�  ,�󆮩s�9��`�'TR�nӚ�����R7��w�t���vʁ��S��NB��R�9�o��XN�W��!����ڪ�{1/R{()�@��̧�C��1�N�F���_s;*薑!��r
1!r�pE���]*񢫺]F����g��p�C��
���ܡ�>12ة��z�A4� ��5�'=m��ֻ�<��;��	I� �iY�dPmdPz���B �ﾹlN�ɞN��j��yW<�T�܃���K�+ �k�A}L���M�*^AEs��ŭ�o �$�Z!�\��[����MzIo�FH7B�	�����p��|�Eze��k�-c��tș�:M����7�AA��.6T��8��K��\r�7AI�(}��)��lA�1�z��31��P��ъ��4S�}�'�^[�
����C<O������$D�zm����7![
��I�����C�;`C�WDz��ɘk�Jm$��R�����e�]W7��k�z�%!o݌)\J�����(&�cN[HzJ�v�%���2��Þ/I,C�L��j}�K&���3�W9��%�怮,h��\R���
���wb�ԍn�5�L�7�;!��K��ײ����.G+��N��s�ѡ-M�j.�.�Ζ松��{�Z�3�)�߽��.�����V_���O,7�L�4��f]��"VwM^�1������/�� d���W�m�bhc�7��YLP��Cm�7;'�^�B	�'u�d�n��"���R���+�,�/�͝��E�tKC��y����lf$?�f�P��9���IY���8������}0�m�<������{�����C�M�-9m�U[��"���.�Y����\|f��m��^u���sy�,.����� &�"�/��a�d���q-Ąq`V���;���������|�!�@�a�X�>I�@��}GF���+�t?�	�z���b#���q9��C�㿾Hzv�>'f"_�p}(��z0\����mq�ŬF�����q��N6T�"�r�HOi
1�"�ŉ�GЃ�|�B��Y�j�$SFT�u4����1ٸ6_b�^�o�v��)�����2�9p%�Lp�h���*�����y� ������EI?�\66����*#����g� �ri�i��4W��D�m�ȼ��m>3��Y��[F$������Lr.�TՂ{ud���G),���rO��ċ��_���*Hԛ '���MM�6Q���{)�m��j�Θ>�4P�з��M�8	)Q$��Ǳ&�k��O����^toN� Z� ��˖�2�/�_�"�P�[�{u�_S����FT�k�C7�MX�٥��f��SL�sjF�����韅6Yz.v�5���.��Mw]LD3�Ώ����vЮ����O^.�^���a-g&�b�nG'C8��v���N��%jH��Z<���5ɴ��o�\�r[Xn�w���KAN����,k=���㰩M�ky��"o������=�x��w���� M�h��ςD]�7m�Y��.�B<d;�E�P��B9+�()����>�p⁡1��N|6��t��§A9y�Ή�G��0-�T�n���Q�U���M �T�n�ޞK+�L�v�K�����>��[�FSs&�K���`�'#}�*&�������8+Ɩ{b��w�j�;��F���/�au<����_M�wR^9�!GK	Ⴚ~�-	M��1C�.!}�Ę[���k]h� �7V����tʼi��=~�fK\������=|J'T#���s�`?�'\��d�8�L�zs�J���\Ux4�[&���`�������}���6�ղu�s	��R���*��KK�_%�+��L���>F�6�͘�����	P�,� Q��A��H�=�8T]�_�Q��u����B��Ī:� �h�0$!W~4�9��4�`;>=��౅�E��!�:%i�'��{�ߩ�/'�6G5��c��P��!�G��>H��<D4CBdS���lq f���?{�M�Ez@����,S��Y,.��O~�TYy��P5�(R�	���i`h #߹�I��ǋ�����v�~�m�O|�́�g��]�H�����5��q⶞��z<����D2�d�;�滈#\s��̕��yu�����W6;C��^�2	?�)$I�����5-+$15�͗���R�T[~q^U�Du)�/�~��]Ki�3�U�*0E�����E�Lh
�٘�� ���xIĔ�Mq�Q�uP΋��������ՆH~0
��΄O8�a����T�SST�8��C m�� 9��`��W��u�����K�~)��*���.�	�H�Y�W���'�.���	� �Ri�[�]�KTp{�0�8���?�Ԋ�#,��|7}�|�����׵h,g/Jw,dK#���Ǎ�a�UǴ-
'D�@Ǥ�0�D�R6#�I�ɋc��%����S���@\���(�[Vf�M�
gN݆9'�ض�>�y[�l�y�8�/�c��KB$%�����%����;ѫl��摍�@D�@keRLs�!Z�GL�����60f��H�� �t�	��8!���D�w
ke��8�-:��֙(b'���AO�Q�:$.끙U��Tt:�d�F#@6���C�Az�5UV����#J4��	RI��r𚄚���`b��9s��'�$iFtÅ��_m�%�`�������v5��iG�䂇\ü�KqD0	�M�������d{(U�q�[���D�#���B {���!�B��!�bqz����(7ؑ�P�"(y,�,�`�L�*�x|�p �CBm���Ry�Ѻ�;�T����*I�Z�8�z@�MtI��Y(����Gn���V��D�NЭ�
��-I�i��ևpB�jgz�E��4�ʘc`!J����T�`����Y�5�?ƣp��V�0���GJ4�N�}zÁ/����IE[��-?j��y�N�:�Y��� ���n�h
v۪�]��Bz�{Oi.��э l��H��A�v��:���MJ'����3ZL~?��O�A(�.�x�"9(��@�ߩC��2�h$�`D�lK�͢�x�X�d�M�ߨ��l��a$k��]�*��jm�O�9o�h6<?=
�û%��N:/q)˸=e:O�L���enL%+^�.���UX	��ID��^�-��cW���JpIk��<��~E��:v��*A�͌+���˺E�ES��R�
��%��~΀c=����jr�¸'w0�V]���W/�b0K���Gز��)^�ħSKx����b�`̂%
�P :y"���R
z��N9�!7ƺ���V/b/ܟ��~s��9���Uo���&y
T����R�� �%M�}6`C\ɜ�2[Q�AJm���2�W��Kƣ��b`i�gGb�gJYט�Y)�1�K�Kw�V<:Y�znP��,"ʡ��P'���]�>���r���G�D���1pD}�y�W�T>�1[��:q�Q� |tNJ�B�.�e���P_;�����:v�!����͘ ��G
���|u`�z�5%�rq�eӱ�X��; |{g��������l$��n�h���oY���Sj|g�s���������h(7)=�eU���e���t�x��#�@.t<Ԃ�d�C#�ʄo�U���A�_AhµC���s��6�{��p����!���&�mD� d�i��(�~]��A#��]� %��J�b�N��6��^�
�t�Ì�H<�)�C�/�5�.��4�3�3}�k�D�Z��7����o5���0���N���@nPѤRςW�s_u<%V
�E6*��S���c����zIdꗑ�����T���c��z0F���&�mK�p���Y?�IbvD�p�-M�&_�a�ᚷJ%�k��v��&W�0l�'-�-&9�B6Qj.[�4�qUWk��'[w�MJ�	֊�h�6Y$�sV�Z��O�"�<����m
A��s�aZJ\���f�I����Z��O��qg$u�i#\]���E]z��L����'�ȬXpW,���%�Yբ�[�u�����j8�\���������E7.~{.�=�线0���?�_Z``��m}9�E�^R/�ä���;U���̮���v�6^	�M�9uߙ|j��:d�A�"0���t^75n睃M�9�1�;̳��+��-Q�k�q�+��=W.��٭��3��I���p��lto$���g�^��Q<m��;�Gk���z_�xEu�s��P���r�z�e���D�Vk%��<V��	ķO��%�����
J�
�ɒ޵--�s�hw�>s����kO�2C���C� i`�5�'Z`?{��g� ��feO��b�y+��mj��[��`�	RF�g��`%����dl�aq��[.G 	ʅ��˃��ղ1ݱO���pu��d��R����f[V̦>��m`��9��R0�I��PQ/d�8�)�$���D8�5RP`���#�L]�r�;��K@��繝Sf�D���'�!�{z�f�����)7��(B�Վ�/Cy��h��"Hr��Wub���18�H6ho��;��PО ������	]� �"&\�Tm"�˶�w�%ψ���$NKr��)
`�;rz#�$����$WI��ʂ�~߇�K������2�s�{��%g�A�h����-A��ݢrf��._�dho���R��Ox��bN�&�?�p.̬N��u���L)Kr~`��>5�� ���9�-n���v�m���2�"C���,S�֪��d�.ɦ�`��z3��.�	��1��o�PY�Y���(��I��`���}��V��K��I�m����E-q�E�oP����nW�Af������J�e���ۍ�|n��D���i2��#]Z�D#F����z
<ۏ|v�����#(=`q�(��DD��wsJ�b�a����|b���#+@C�fH��b�z1ob��-���{,�����<�2��[�+f�e�*���U��R1I@�߆���l[$�q�n�;M�^��z��hG�eW�5XdX�B?ם�R��Oҙ���&�h���+��2Yq�yU�R��x�21�(�GB�|�m==}����9��1˭�zs���Y�r�҃U���Ԯd���NЍ�G��|8����F����L��`�+���^�x�q�y�>�*�&*��r��k�h1�<�b��{����g����>]s��oA-{L�E.�H{e�v憝T�7���'X��P?���`�f�V��a�`�B+cH�D�8�K�B�����X����і��0�=�m��⍤��&��>�7�a��	�����$��E^@_��{-�e� ��d~���Kp1J�,�7Ң��C4
~�ɘ�>���ESq�쉪%v��}
�����]��맞�s��fTnROǊh?_ ���.�@0���y�B�Nي�s���8%[��۱N��FS��.L��i�|1<�P��?'@�|�� ��G������#0Rv�R�9��J"_��G�^���N�>�ԭR���9��l�����Ŏ�q��7�Tcs�E�{�+��F��ݓ��uh*̖�; ����4̋R^(�О$�hx�����JM���6A	���e�6�{#e<��6���w���*�f� Jw�M�x>��dl>�X�����ڲdXx$���-��l^J@]�ш�����r'ó����!��n�WX�R�b�Lz�����������Ӫh<I�CF�.�=�L��mP��B����Z,>&йᎦZ���;�~8�!9�~8��_��s|bZ�<u��W~z&;�5�ɓj["�C��U��$y��;��VR�c�ÔyW�{�1�i�{Q6���	9P�v�>�N�W�\��	�򿸆.|�`k�-���e�=Θ}�C�^���YBg��_�L~�8�7��דsm-L��܍�����>(�|<A�[s��Nl..�}�V����f̶��)$D���ƵPtl�w\|��C^���µ]�Y��K*��Х��p��b��3����\4_T��aX�	�q[�rCŴ�����G��Y��x�*d\��
:Q����2�"��!�Dy��hߒ�8�bq@t�xH���ίmt�F���m}�4��8}���U�5>����g�%	Oi�;�A���i����V8f����fj�՚�DU�����6@I-k�W��S���=&xt��o��]�QT�h,"9=!��~��\l�t��ʜCiKO�#4.�v/Ru��s����Ro�l����"�r��	���[~]�"�n�{�r@$l/ʻN��O�.CȌ��n�HkLOT ����3��1�ִ�7�)F0p�ǌ�֓��wۯ ��'pSE��R@W&������9�Lr��+��.K��9s�V�i�~j��AET��C��dd���T�{�K��A6�}μ��;xp�G9�>~��8H;_J#��|X8�Rh���e����	˯V�_H����dv���Z����M�p����g=דQZ:[/q�dVS�N�zC >\��y�SyG�� �P����8@d��B���A��$�k�kt��rВ��kd?NY
�v'�l#1��A�]�^�����kβ�(w%&J½��r{�c �A�u�}�H#`�L�(�Z�F���r<&L��<�qų�|�0F3l���1�Z�ђ���:���&h��h����I㐢!AN��ϻ�ޑ�̭Gh�����AZ*�
8
3�i������'[�e�������A���4�9��q�2�t�7`Ft�5�L��;� 촏2�|���oz��n�b��jؓ�:�4�{k���iBG	&��%�M���{��и˭]x"b�C1L�+�����`�@�-d��z���SU���+���l����i|,S~I�EB>d딭u(WR9څ����K���M� e������]8e���|�3,��nӱ����z󶊌	z�S���$M��ԣ���a�=��*NU�:��w�K���jx ~@>�6��#���
����\R_8�[��ߙ%tC�w?ʹQn�l�c��]1�:�~�v)ejY
�v:/FXHI�!�Ķ4�UJfٮӘ�%���5*AW�.�n�ߍju�>t��M��~h���n4	e�oA�^aB����� ��1��'_��p�L)C��O`u@=1ݏ�fѧB�o���E6�T61�=R�����I}�%���֍��s<��߄��f#��*~�W��Ėe|Tx]�����7�P�p�yc_�G�M#B�5|+%����BD\��e�J�/�º!��,��?�%���<���6��#�מ��w솹g�m���`y�1k}�pn�zVAg[��Ӷ�E0��� 
�}���\*�ڴDs����
ߐ�v�>w(��ڊ�1kT9���p81��ӡ�r��I3�	H�/�)8NV��
 ��7��q�}�����b%�x$��D#�~�;��q ��Z@�{R���`�Y�ȅ9�{Q[�����g!p� �����t1���7f�I�33$��甓�j�X�oc�E��
M �,�K���ao��`6���h���-�����ݓyD��������]���'"��w�&�6'�E|w!�D��H�^hˎ�� ��į͏���au���	��9��su�n������ Y�@},��?��x���^RXб��Oerdk�oßC���J�|�yaa�v�8�}���z�1�'�wnq"6� 7Ж�]��֐��L�+�A��G���bZII�q](π9�a�z���e���T�UR���NV��d�@ki�������$,��k��kЯ������FL��;�+M�u'=����q�����6�|Hp�6J���Ǟ��t���MCs�ܢ;E�}��u�O����m3�z���L	�Bg�@�}�u��	���jǪ��S�t��N��a�;���T�CD�+P�v�H����Db��@MἷQ�o2�ʜ�u�8�MD: �>����(�����gY^HM�e���NH,Ca�]���Gc⃜��m"��F�~�s�������қ�X���<�\�?�\����^p�J�o��z���zg1��)+���L��#cV})��yb^��ƍ�U��g���hc�|JE��B�0uϪ�(��'����W-���΅u�M^�db��-4&}��wz���2���ێ�ȥG/N���S�B<{۪ ���f�k�d!O��_�]��>�ͅq&ɗ�)>�j)�ku����{��L-G��q�ⓟ�)b��K���x�~,$O)B5��@l��]
z����̟���B��4�L�^�P��"1��e�{��$�ܟZx8�zz%�ZH�Mt=Z����b8�i�xJ��?z�ƫ�jɁ[Ji}��`b�b�d5.����&��t�Ek{6�����Ш�_zd�����a������QC���Ӛ�}�dmebt�O��v-�K��F���#@yx����`F�C-0 _b��?�[�hF-H�Hi��r��vrtFd�����F��s���ǦUw�W/�&�x�ͺ�M���q��k�(k�>�]+oVﯛC9E��#2����#K�Q�L'%���`	W�Թ��1t�m+Aކ�Z�w_��ք�[v�F'Z@�������c;�����q��t虼�=�ـ^�Mw�/�C6s����u�eL~�쎌�W H'� >e�L.��}��׎h!m��!�~lbQ��~I|��Pj	���S7֣ߩ��X�6�ڌt�cMz-UԻ�7��Yp�"��;��7QG��=�Zq�	�yz�9�h9��i>A�9l�X%l�MLT�c~MR9>Oj�	y����PKX�6?��f��[P& �6?��Af�}��\ҡ���28F��Ж�����Ꙧ����`5�A��k%F�\8�ԉ��vf
YvDh�������|A���F&G���;� �`�b����go��F��s&k�ˎ���Ӕ��+�5�i�%��g�׉�	;KLZ�Yf�ŷ��-���!rq��x�*�[1�A��?W`��)�{���MQ���<��"�6H)����1R�$�e�9�g�Lι�,�����ͤۅ���Y��0Q�Naf
Xٟ!(����]-b���]A��̢nŪ����%_-���������/!T�7�Ui/�#wpZ��&�t[�&��=3'r&O��.9�7�aM2�V��5�[I����/�?���@ij7a&l���*�\Z9�]<�(����30x�3�~]u�U5;�UY�}X���?��e��f�|/D��D؂@Fo�ߒ�bb��ߜQ� Dd��ʺ�^�=���h�%c�������v?�rw�j����D	k�A~B�!���k��G�pi�4�F�e��O$5^��O�z_�C��6 ��]�wJw�&�A��x�{�Q�G���?sq�>Gb�S��T��"c�(jDqu)�ɫ�j=�C�w��k-JlZ��V�bI�#[@�r��ؗMk��������A�+����l���t6��Gy�<2~�V�n�G���XWNc���'n����7pμN���c���~�6���%���tT�P��E��@�d8�S3[�7�6-�:�h��oԨ��|��,�, Ĵ���Vo�C��� S[�jOGH�S�u�b+Nzʉ�h��u�o�������MF$@Ѫ��aa�fKL�t�$�Vk ��Y�~E|���7
��v�6|$� Ȕ{�Ɔ��ѱj�H3��\jͭA�T+�<�xR�Hy�3q��!���h[�xA�9�˰Wg���f�"S�A[˳銋�n��y�U}�E�2;�̺#�V`��vÃe����'7�Kv9���	�ð�fd�
�F'(��\�ߴ-�7�6}�y.�Ŕ�����mRL,�m�M0�۸���f�ǩ2���)�˙΢�#6#I ������wl�?!5��׳������K������A������U���
��v�"cH���Jd[Z#����`&O�ǡ����!V�~9A�a2�I��WH� �9����kEQ�S	�s����%��uN����ƽB{�BX�;>�����Q�U�Mk��	rPc�lO����Z����&΄T�%v���h	Fp�D����1P�\�"W�X ��X�_}��ԥc(84�9.DRb�h����._[��J�Uv?Xuy�dQ5-G���9H���d��5�`�}b�T��FI����w��ʞv�+@c�|��$�>>��Nk鳑E7���fk�D��V���}E�A��1��T>dx�ɛ�QS)�I����0W�`�%�Ӡd
r��4|V�αn&:��]��Q-s/
I���(7S�@�f2�\����N���P՞KO���(�Lh�����A:Վ���i}���&���l��:��:��k� �"v���lD��y����W�#_W��[�8�����C���<�4㐨B\�G��p��g*W�c�k�I;8�� �/I~/�*��R�n�Kr�y'�d��I@5c�')69�R�T����L�������
`�!a둠�@�a8Z1Ԕ��D�>߆����^�;�i�B}ׯt������f�����K�(�D� ،�hºY����}pT�Xs�����+{y�J�W�+8�;�,7~a�U�8�I��"�H��@4�x�� ����>~�	�'%��<yB)ᄻi�,2�]e��+۷�+"J:g8�/�}��`��(߆͉��"�L�CQݛ��$�nK���*O��rR�H��fC�18�m͇%
�_�Wk�a���v6�Nf$����P���U���T�O/nQ�H��SD�%��_m�()ny�A�`�rX-6Ǧ�Xhc��4̹�*7Y��k_(��O�z�S*'A*p�|��v�kg��J���@M�����������3 U��\���xȆ4ƚ��������k��չ�}}[/�AAW�@�ڽ��}�w���}#�<K.���� h*E�m�&:l�!�,+��7��8�CO��F%zC��/�y�|Vj~��fn2'����X1_���gs|q���jEI��A����&�����q�[�\y;3���:дD����P�<@��t�S֬d��ga�Q1N�9nor@M�&u~[b��P����|�NL�����EwkUD��f�Z�9��W2 ��0�ն�ש�d^+����1|�k���{��^B�f�cg&RץY�j�ӂ�ޤ{���VPilG[w��u��<k��6��q+�"��C�����cͫx�[ ��EA�`����Q��a y�þ����P�g_:6υ/���~,��`
���zq�����5�<�` ��>d��L5�3K�oɜlp�%-N�-�;w�=�e�3\um-�A�|�'�Ҡ�x�P���)�5ơ7.�K�o$D�vKó��L\i͛��|$�n5���9���[��R�&?F*��:��A��wJ��I�k��Z��%q��U�\�2�E�$@�cI��>�^w\�Hb%�\n�-��Q!c�ܥG����!X9�e�?k�O$��B"��ԓo�	W߬��e��eĶf��*7y׆���ܺ�R�^�<��! �"QX�&�^�܄�3��F�r�����!Q��HW�n<�&ΏV���k����HV]PMx���R��	җ��+�ﴭ������%�arp~<݂���S�����Z�F�έ;�5�������t�)ٱ뙑QpYq��U��,�!�\�jl�!��q+ ��+������R�L��i��M6���ݜ�h����j,�b|��y��l�+P"�bCE�k��ᦛ���9�v	.��Ͷ~�d������
&����������}���gD������R�˩��.�_�)�,�go�Ne���U}z��DQ�@C�@V������� B�DF��c�i(�o ��(V0�v�V1I-Z�G�N؝�T!Q1��bT������Q��Mَ�֗���os%��?'�K?�����B����7�^�7����3/�M.����ˉ̼�LT[�@~� �P4[����6��t�(���:6Z�S�)��*T#t19&铔?-�a�#���k؊�H�|�6�L��$yZ�RTB�+j��G!'�ڟ��:��op�l�����4o�2�{�.k�z�������ӹ�|z[�lb{ȁ����פTUo	�v�}̐w
G��j.��K��ˋ���+U�ԏ��0dy&�Eٯ_��h[:��NgrX�J��k�hq7�^�Hh+A�OB���Q�2=&[,N;�%����]^���s⺻p׼��(�6�_��]�c=5.���+�V�ځ�M�j�ٌ����s�.�y�g(v�b�NL�+z5u��e��� ]�:r&�l_v4ҕ��Г� �g�3�- +NG���e�2_J�����^�@��u-�}��D��Y���"&��+��A2�4���C�
��2�CskD�k�]]��F����`��4��{'A�o6tk�aU���l�7zD�T:d���a�;Ý�z������S�I����ֲI�1I'��j-\�S��='l��U"$�f�#rm��ȍF'^b��.R�?LY?�-M�粠�b�x��62�ңS��!�5M&j#�� ܲ)
��7����v�Y>\��sc&NB�Z���^vMNz��>*4�j�l�Ε�d����d����B-A��o#�,�l_N��($�!�������2�4ˇ� �Pρ��פ����Dj�C�b�V��[�Ф�A�ٌҳ�To&k�?�/�ep�z�|9H��ʩ&5
zX�Z���f~�xz�9�e�j�M�KP.(ަ,�Q���w59�+�c����*��FS�h�3Y�.��ʡ�>�o�X̿��x�N�����Fy+���}x�7\'���zg闌4��L n���G��y�)���Н�����qh��:�������w����E�>���Ӥ��W��u�x�8M�9~?���� m�"-�Bx��1�
�?$jZ��0��]�yT�A:�(�ؙJ����?<'���ޜ�L!*�p�Z�y�ʘ�-� ������Qq��-�i���s�1�Z��(dZP��C��N��>���p��@�����Ǥ����	�h�z�ܼ�����t��Txe�cX�6�g4#a��)��Ȍ8Y�v�Ǻ�ϼۊ�?�.�Q�.z�q�����a�Yh�K��-���Te�����$Ԍ�f`�w�S	�(c���|��b����`�f�y��R�������a�R�.�H��V�.��QS?l+�U�#U`��Q��	1cP���<�Tg�a7 @��Ir�~�g���>����mB;[����Z)f���ǋg��y8�z��m;�K��P�LҜ��F�5G���i�9g,�/H�t�Ϟ�q�6w@�f��R�T��l[��8&;�"���D�{�[И�L褏��a@F��D�J|��egR�H8;�-��ǘ����C�K� �xU�S�
,���Y~�}%G��g�Eka>��_/e^�.�bt*f�� }=̼.�l�7��Z*})�Y��������/?g�#�1D��a;jΆ�a�U��G�������L��Mᡓ�/�Oֵ��~�l��)�9��+I#j��&���1�e��K0b �7~�Uk!:8w�]/;�)Vg�o��M'S�<e4sC��vV�iV�;^V}�j����/Z���2L��Ɛ����<�N���C�ߡQ?��!(�z�k�r�=\Ś`焬K$�Oe�Ʀ�� ^��� ̃�\�?�aP��0�fR"S#X�@
վ���	�����}u6fK�{(�i�R虷�Z���a��"ڨ��N���i���׆�{8�]�Xr���yE�!o��? t�h��D����O��᧚PV��WQ?pC�:� 6��.�;�T$9�O'�^�3i6p4��|� ��oR������5z��B�[/:�q�Vz�/k����2oWeVZ��J�\QpT�WkN.�U/+�����8W������l�>�&��#7��~C�o����k�:9�_�/��Xm�O�t�Av*ģ�#�0?�il���W�j�V]��Vpb�,8�U�9��~d0���
3@kS)'( ̘�=:���
�q"�^:4������Β@],d���	�t0�=�U��ol��@��t�[�a�s����H�NBL�~r@���M�S�Ů �F���{H�� 0�kd�g�<d���^3� l����f�T�N��(u�n-��T�k;���۴w-���8q#X�����.�������ZS.{�=����f�yrM}w�'��ˣV�o�b$���K��޲BZF�����o����X�Y�_-:�N��d�Y�P��+.�5p�U�\;"v����Mrs�t�e�M`��3"�:��!�Z[��Q�8�E�1x��|H�.���yW��>�9�dI������O_� ����r*��(?KBgݧ�̮��_1	�d����΀eT�
�r������)/Go�z�4sL�.���E"��ߊ����qU����B�:�Qya��Z��Q�kF��P����=�+z�h����97�$*9���3K��f�wO�=_�t7�z)Էn��"8��+Q�\L&؅�"�wދ�C�]�L��iՖ�Ɯ��I�Ix��XvG��/�S"��t�N�;H��g��"�I�޽¿8�/72����A�� �c��.8o��#�B_�qv������9n��?�,��&`n��c)x�U,Ud�qgUP�Z~V�cy���d-n\)w�]����*�*�ww8�~�+�J��kk�vKWOd�ӛ�[a,2��I�NeC�V[c�����i��NQ��6�$�����_N��%��c�)Dg��|����Z2p�<�A����r�4�5��\��^v�c۩���V|c�`9��+�P�L#d�]���a�T���M�z�Ί��m��qSM�~���r������18,��\
����Z@�_��fc�:��4^�}�s�t����q��S
�D��	�E6~�=@})����C�g�aQ�2��`�������I�6�۟+�$Boo�~��Dl�ȪY!!z��X5�>3\��i�h�6tCB�73��~��N� �1ަ���.��,좐曪s�S�h�6Z��|��:��}gs��!�ٴ�p|y�E�o�G[3rEi�+0�d�jgEhF��C��՜��G�'K��E�O�S�ss�kЯ����+v.c��@���fc����M����A;B�L�G��� *Op"����1��0���p�Y�Vg� Q*$���5�E����+SU�}�Q�%'�I��Ty*��B9��h{*�9���ƭ"6<F�܊̤ׅ�OXN��S>8���ֳ��f�@�����!��-ě��Z�iP�,J@�����{J���E	��5_�w�������V���j�B$ף��Fq:�V���љVjb���,��?#�a��j	�>^��i_��C�����G���yx3��z(h�q�CgG�� �����D��
�ų������l�W�1��<�Rב}%�j@�R���K����<�"Hwb��8�#�E���Ô_d%I]���3őD!�W�n��6�ٝ�7����)q�`����>�+A;{6P��'�x��e=��H$O[I�cZ��|dDID��p + 1[a��b�C�%=1��g���H���J��UAV3�nl8}�g`r����u֭�s��<!%�ZXo���G/Å�sә��q�(����{�C��sM���\6���jvI�ւ�6F���e k�W���\�|V��`ﱐ�S���y��������麯g��N��W�,ǘHnk&Y�W�3�\/�M�y����#j�#��F�G�5�z���[�����<�s�Kb�(�r�~�#['�#��\f�ʔ�u$0'.�E�2.��nB[a<4#�a��@�?���慕�w[�!�ܿ7ȷ����G��8iX�W	&��K�[sM��Cu:�9q�!��N�����`{�y���ϯ�]<0�7��n��N�v�&#W%��H��W*bw^IUsK=n?��1[������K��30��T4����E��c]��)�>".Lj�!�e�et���{�Rm+ڨ���z��Yl4�� V�S���Z;vq�E}Xq���$��N���b鷋GK��D抙��`�0���T���F����\�r�K�a��^�\8��#�YY����ޤ�l >J��܂0�v�)�?���,Di�˾��@/R
���:��u�}�Z�z���ٹg]��:SQ)t!���C��tcW�>z,���(f�$�58y�"x�e`�Z-����50%��qVr笐����Q���ֹY�m�����wm�؈�?b�!*��`}��bF��]��1Ĳ禮|�X!�� F��y��)�����٥Ơ��c"Z�	�fkp����¾~���`��u�!3����\��`�F�L�MwiẾ�g�Sf���jO�;��Y�ʝ��`��"�@~���V��5���T��Ms�b�L@�6��)U{��.$b7q~u�.D��H�z͡������U
���:���~γ'6���?��⯋h��`0yb��fs7HE�1�ЪX���X�viH��D��=˶�	���w{�P��6�Ƴ�t�:K��k��Vu�+k��\D�܏�~y�rn�TC�yD>��4�M9r��9RW^$�F��ˋυ5�`N�N���)��>K$E"���_�/�<�$���k�r�!�Ǐ,AM5���j��"ΥԪ�V�Jj�RZ�J����_	-��$��}���Dac/N�O'����*��� Ӻ]�0�B9���Ut��	�7�U{Ӕc��9�̢�}<��#�wCK�i��Fy��)iD.�Ja�>��,������E�YN�'��
�R˛����dBɌZ�՚{`+Sґ��@����d3�$�hUla� p��lk��	�Ĝ�ވ��	�*�5�VԖ�$oo͖�/'+�&t�e��s�"��с7NP��D�X�,w����D^���_x���	^\0z�`]�u��0��u�I�U�A*iy~�%\���^9��z���yL�C�8��獰����K��.���x������ď���\I��2#X�t�%�W���h��e��c��Y����`�������S�
z�t�1�0s͌�*n~�j���4t��VwН l�u�ޟ�=�����֏��7���J��Si���j�<�q��Y\��u��=��嫜�����3��LV���� !�y�||G��*�D<�|Sq�N���'w41nl��qk�����9c�`��A�$G���E8���h��xx8ˏz�"�o��ܕ�_�S *���rA���O�(�����q2x0��H~ǽ������7���':/^�r�W�Q�'��a�GR�*ϳo�����<y"��-�K.�GX��Jq~e��s�jH���,��N�٥���:�^`�d�GԜ^�/�Ь�z$X'��o%���i_�n���G�<�Jp���8�k�Qb�P|qV���mPYN���4fټS�U7���ٓ�ڭz�t�jU����58� �L��אG��MQ,J��;�&�M�5�6H��
��H������35=�".{�vZ���6J#�;|�v:"�zЄ�ä2A��	�wBRXѵ�ӟ�6V�/��#ʞ���,"\u��hK�ׯ�CLc�c���-ԫ�w
;D���D@4}�����6�-�����b_m���]� +y-�x�Q��UjN�d�A���pqSf=K�#k/�v��l7e	`l»� ��uFvWy�����9<��j��AV���pq���sYh��V�&�:�	��zL����t�lY8���s�.C.[mǀzb��P.�,�o���Nx��A���@��M�7���Q��e�r	�\�5z�7�� F�����F�č�bV���4���'Yuw��Y�*p��fЏ���EB�T10%�d'�[^�k�	�c�$��7s$��abI���f�G�JDM�+7Ƀ�.�F�"��X�Azx�	̓�n�O�R97UL�(J{����u�>/1~
�7]��/�8�ƥ�l���C\%�䤕���y@�Y����Cx�ܢ�^�v�"T<�oz5��N(�UY����c�oL��h7j�������J/m�ї;dd�ɚR�߸'lL�V��C���0�#m����?�f����v?s"��!ʄ�|�9{�+�R��7'��.�'<k:���G�gi	���t�(����.�J�sѻsR��%F���sii4/ϮO/_��]�T������h��Ո�J�cٙ����ū�R�W]�p��4_׮�~���g���K�rM2�
+������(R��h��*-I�Rn����Ǚ5(�q�ux�������3�h�!�A3m| ��CM�]��闡�/�� ��������L�l\v�fr$d�Y�wK���˻mC�=�g/���!����V��|�q1�|�X�j�KOkޡ�
��l�	��[�W��g��!��M���񸑃�O�������M��ٸ�����M�б!�����:%�q�>�����2�yH7�>M
�N�ѭ����9��!�|��� �|��<8���b�à��&P`�ۻBf��4��k=y��ȾB$����hU����P���ٔ��?��x�H<=���!�t&�U.��B��#_ ;z�8/�����j�->Q���˖U�ssT�'�EQ��9���e�Jo6�:�pD�@�+E�͓o�vX�~g�d�4V�(�"Lp���X�d��,.%�4���_.E�&�7������l[]����E����*u">)fՠ�ߗ2m	����B�q��PV'�ÈWMH>�⫔��8���m�s��q����.6e-|�|F�*��\r��k�V�ul�vrK���cq^&;&�c�T� ����{e,Eey+��|!������p�����q�0/;h���9s�㷪���y�q�od�e��A�Ǡ�J�ed�����Ԇ�9
��V�H&%� ��4HM.����f1[\��:�w�V��1&��xmE��4J��t#qǊ3�n�-��ʱLI�fr��5/!�y"讨�@�Ma�/�Q�n�	VB�%�i&�~s��M�������}��o���f��B�$��y�+mVtl.P9ڻL�)�C�V~ȼ��\�b����\�Y�g���r�`+�.m��
iR7�ث�s����rO��C�z� l�1������6��K"7����&k1�)Ɩ�:A˯_`��JUg�nk�01��NS���Ͽ�(&l����C�x�0�=��F0̃�e�F��W��&�O;��V^�;��9;�Q�����[7�E�Q�!�|���t��}n:��-�5���C}d�L�;�Ñ$|��m�eE�@��а8�Xvc�I�تf�a~���˹��Pޑ��M�@�(l�뫩OZ2N�͂�z�x^mը,��}L�S��+�g��_��-ً�>�B���B�F����à�����C,���Mp������gȍ����Nq��  l�ܐ�2SZL�����ֿc�fO�#��U<+������Ǡ+�M�ɖ�`"@�aE�d�)5#���ĈBu'��=�a�JK�W�V�*cV"Z�|�jZHI������D8��4C�!=�Ր���5�����8>�֓�s�b��?�81���l��PZrЫ?Ɂ����9�7�i������3��-rp|�	|s���?�Yť���]�R�b�3`��H [���7e-��E�B�a�(J�A�����F�}J�zQ�#��o]�G��`�;��N�R��)������-tL=vAH&�ᙛ�k��\r'�'���qhUd~͝X	\��MA��Ɗ1u�����KB�$�Xu�d�6�FW�o���㉁������o��'�c=&#��(�����-�{�%�xFy#`�EFf-�B��[y�?�>����DgzY*��1j��H��D?��'7r�󙝬�}�
���1)x�Sk!���R���%h���,�q��¡�Y�+�ǐK�/��F2�#��y��c�}��~���}�(jR�Ί�ۃ��r<������	!�5-s��
f�K���@�V e\�2F�T�h�Jz|T]^JA�1��a4Z�ھI7����?���_�.�[F�7]�HS���qrci�N�ȏ��m����05*me>��&�vT�v��,���)����)�)1tb��1>KTT��ee�R�P��-��� ٧%�\_����!�2w���4`R���O�U�!�σ��Ѫk�]z���b3O'�W����&��šE��ii�������}���?'�X��nU淓f��L;.���{����@Me���S���-~tV��e�D�%�׽{�� �.z����9Lx�P�e1��aZ��#f�(���� Kđ��O���+�t��G+��u�m����`Jq�T?��hq>UP�8�V�A�yvd�y�S���ÆM��9�5����nC&A�}��;n�'S�ʯ�r�d�Z9��A�:j8�	�� ��doq��L4��� �����h�A�l3�9��tr���v��#�p:��/&��p$J���Ј+��˸f�Z<>��ԕs���˰��ژ��JA�?2�����5�F �`��� 貟ګ��"�"( />W�>��W�\!`�7��٦%�NG�cρ�@x���ז��H'h�������@�(����"�y�IL�!�v���5�0���W˺��B/�D�,�,���y�F���n�(#W�aV��5�?��Jg�~h�o_���� �:�R�1�i�R�+����C޸4��a�oJq�H6X��F�H.����@ï�戲(�4��AIY���dY@Ei���ŲS�:�D�Ȩ��iX|{V��p;�p�����eB\�!�	"�=G:��"�c/F���1���6�����p˙�i��|X�`Ӣ��Tʶ>q���r��v�p�\^�Z>��5{W�|s�k棠�����=��T�QW���-	+���}q?S>��q�x9�;MB�=З|�s�l(���l����x����l������+�r��stx2dc�����d�uBl���)6��n����L��M@�U~�ySv�e z[� Q��
��h=���F��W������ps�#
��:Hx'b�azm�����$�Ud�N�H$X&<NS�m�.+��.�X��F��Q����_���mT�n��/~�7�in�ʳ C��ߣ�_�Mn�9-1�%�gI�o����"�T����ӲC����&8�ц���UE� �K�4�R0�oju&��ܙT�c�hP��~
�_} y؃syc?�5b��6=
^7�,>hy5�(�y	�m�x�`�����u�	g4	x�*ևH�4�!-X�����.e@��2��-��(D�dӶ�/�<"$̡eDk�G�B �f�5�"����g�-�E��
{���G��y���_kĕ��&�y�l�i�������N%Aw�4�T��~�YLN�-ׁp@�doO�/���Vr���A��>���8x�.�I��k@Ⱥ9���%Sۺ'��gJc�}�#q�JW�yfiK#��ƶX%ز��I������S�d�O�bDpI�r�� �1z���@Rv ��8Fq�ƨ3h'����j�M���O.���<��k�M�~��P��Y\-���HK󔿉{��0���ĳ=�&ֆ�W�;�Y�' ��`���4��Ԋ�5���s�Kk�1$�/
'���:���Ƭr�40����N�6�ƙ(�z�n�p���C+�A��I="H�x�`������,y���G
H4BVVP~#�2m��(���.���6׀Y�XwPW�}�����Ss����*�Q�M\�)��@$؉:�륾��L������VJ!h&^��y��6��,��+r���TT,?h{A����hċ6XA�δn]=��k{� 	enϪ��MѩT�.�=۞B�|:vK��zGo���[3���*�lZY?�|F�T-�bZ"
|�ŲOy�)(��h�W2_N��O飯�d��c#.����r�l]>�����e��4i�����|gG���~�p	j�J��A]���~�����Z5n�"	DZ�獘�9m�`~҈	ͽ˝ф�� &�A��
�v�h�x�a6?�[�[�cBa�k"�7��:g=&�.���0޲��L$�K����Lw���[�݁�w�K�,n-� �,�,�ɾ �K3��
ɬo��lgs�63�������Թ��
I���s�ҰbS�\p���C �b��/=g@��Ѷ�A�+�j��ƭ���=Ts�n�l5����:�]`#X��dϣ����x�8r�� �I��Xy'k�L�%��29������+����қ�o�W����P�������t�̏�=�ɖu���Jme<%�q�i�{����G�H�m2���$u���d���:�g+�\y�/�����VX>�+�t0��X˧�S&��9�o�Fw7�}W��J�dd���nd���5u��;�"�o���[o�p��,	d��W�I��>#ll�L�F^�euV�7�9���5��3����1/g�4v8q��nByB��q��y�"ʧ�#��71�#��<�u���c�ē!B̷��8CЌq�㎆��.����d��2�r�1�s6`�e'(��j�Wy!~�J�/�N1�+��w��m~��d�Ԉ[K����*�W�v
7E��@p\�BՁ馅�4f/�d�*��m����9���LD؁�X�@gڎ�6 B`���qbk����E�?�y�{�斊�O��$�T�ʡ�8nn� ����ܐ��W%��,'�5S�dB�e��	�p��^Iq�Gun,�7��{��I*�z�M%t�C0G�4AW;*�)� �����9�Ǘ��w(�mJzF�y<�Vu쯛�AgYo�
Tb���Ds��^ӫ��#^���u�i?"�x�k��􇀀�����K�D�52Ob-u���sr��'s[H��:���'�p����b�qh����ڡ,&�|��6�����9ы�@�OO�g�I}zLPK��T�u���g�;�s��A�{�Ƶ�|���K��-���RpkA^8Et���da�LH̥E��K�<ڃҠ������0Ҁ��b8���o�mu_xȇ����A�HqW��Qy	���":�RZ��o1>`��  _x-��g\CNvy��Y�m�ȩ��#��D	3���J{���S��W����:j z����Q>�����:W��N�Ñ��>�$�����.�h��ZQx���J�>�?-���/4�R
��!(��|��ł���v����퉢�XY�[2	y��������L��&3���|�}�O�;�{���������B
�<��c�n9il{��-���}w��d�ʭ�Kڦ�����d[n�:0�z��.:{zH��]��woG��JF�scm�L�"
Q��E����v��{8����Ϣ���z�~xӛe��n�&��:?����D,%dUl;^S�A]�|�����������jYa�ɒ��(��v� K���|��U��G~����I�DP���>w����tm/�-Z� 
p�����-u�=⢀�Y,H7P�i�Nu�2܋�a&���e�7F��7!\[�<i��_읽	�H�^(�U����W�9��ұ�>�ֶ5��\������$61 GqҦ��Xj�qs�����}��s
/M^[����Z�o9%�~S�5�\z��K��m�c���X7Q{^?�$�h��a�&��ʞ?��:�D�#�Wٽ>J^�wX;�cpX�톔�pj���8A���+3�ϗ$ �Q��%} ���Oy	.��`�C���s�c�Lx/����N�@}���"�˻�1�(÷ō��8Ä��&]�9�"���x�6�/_j?�N%�k��"pu#.����U�L��B���2�;�������}��1�Æ�0��8�Hv��	�%���#"�%ml������V��bC�1�%� �P�?�חk�'�qhD�/Kr���|%4�j2n�V�ĩ�b��k}X\;�"x�;�z�����e j/C��ae����y_l��o#�=��!�DSi",� ��/�����Zvi�~��B�ҼwD����uC��lI�9���蒏H�r�ա49�,$�� "`Ϧ�ⓐ���[��%c���$���^#��j�2�{j��Ӫ�Um{��6G�@��Vd}�@�Ήo�6������:_+ƾΌ߁�]􈥽�ozK�F��yQK�|SL�o�]+� ��8܏�N����23q`| N�!��*<X����7��#�12���	C��[���{ �� ��;	e#>p�����&k8U���є���}�_W��fU�EF�d�Há�oвz�w�Ҍ����Kk��5�.*۶�nd�,�a��R(^�/���P�U|Y���N憙�0h�G��n����t�_k��L ��$ .O:xr���à�B\N�lM9ތ�CXu��K{�3% �}�!M��ҌP��vU�,A�/�Z����
�?eȻ�̚t�� ���b<�0]�C������-nuWt�QOzLW���7n��DR�eE�	��l�!�!�i��W��2�S����*���%��ۘʞ������.��r!��|*ߧ����]��^�y��OE�ޛ��W�F�/,��1�#�����,�	+z�w�K*��Y�_�^u!�BƄnP������v��)��"~K�ɩ��ޒ�Q%��.;<�<- ^�p}*���H�ŴQ�m\���`��=Ȇ,� ���`[�!�%��vP|�a�|����.�wΞ��F�֊oF]�Z�)I��`�}zo�߫K��Tv��$x^wO� *+�x�!�T�p��9p=`�d,����-ȼsmg>��i9�?�H�Wk���2�ZB0]�QS"��uSh?o���>��Ċ���]�o���M��3���Q.�42n�n��r^L�f��f���+�xEEv*�Hg���]�kl��n?eP����1���z���H~1���i�3�v��k{M�1�pz)�M7w��!s��w6����F�}���2��H�E� ��"���!���k܅65�+��74_)p�['#�<>	Yy@x9��t};ce�u���0׍�X�'�������(Av��p��/w=
��ENҁ���aa�0���+]o��%�_��QE��Y�Ӟ���N��B�T�0=�zI�S��8�[���é�*%~?��Y���S�N9�@���TV,���N`�O�ר��R�G�b�џ�Y9s��xV̆r�[�NnSv��s�$�D��G,T��eJJ�z�u!n罼<�VC���`���{�j��k$�������f^�"�T��0e�¦�[?!���-\�52��`j�b��8ԫ����o�,'�����?3Z�>/:�nq�|O�A��9ܽ�k	��u4QO�({�l�f��c#��C���+�H�k�9�\���xQb�W.)�KU�6o9=)pt��bӸr��g7V��y�
q�(�|thP�G�q��5��ء�|���R�˨����zMZ��~� Rŏ)�li~�8L_�q�����)���ḩ�9y��!on�8E|x�°��ǎ�Xk�1ȜN�[��:c/�ck2s_k��s:*P�%0�Y��B��X�F�/d�_,�N�-��xw]:�H#s���;��r�I[�4:�� ��D�je/��,нl��A��`va(��N��8�|�nW"Zp9;���~��	A82�H��F�:̓�a��c�S��~aD������tQ�\i3�Au��e��%�9�(9����=�H���
X���7�t���,)�O@ۂiJ�y%2���Q�'7����d]��V���?Sm�G�0�?Nkq��!��r���9c�Q �޲(�m�7��DPZ��I�������F5�=���صy4����d�ܠu(��^O��~��@�.wS�����,�f���7n��;kxE���c���}D���'4�
���U�o��o57�[g+�@.z�T���
��N���Xh\����f�Nb\!���@Q��/�!"rjL�ξ�"������Rd=�LC$����?�ڨ�m�y�*ԳɈؖ�>Ñ<���(�|B���ALF~/�ǖz[o텙��߀�ߊ�~�dg<��o��#��4�������yO�����F��7�;�Q��P�ko�g+���.bw�⇩%�cxn���V�'�_���b�G�Ǽ�}�5�f�(k�촏:)04#1��ߦh��vd���:������5[�'��D�C�n]�^�pR���i}U/�X�	w3S6ݵ� �=��0�b�R�R��=:�`��w��������8ߓ��m�k�y�C��+���ھz�f\6�

�<1Ou�u�M���E�s��&0Q�G�f�<*dᩗǫ�_�ٵq喳�<�b,O���@�G�Uq 
:�o����aO��0�M,뺨�)��_^�qզh��
2����aF����_n�|w��hũ1Z�o|/+E��:��`�+1��tZ�j�%�Aa�ᤉ�g��MW�k}��GQ*%��X�[ta�Gʫ�q��};�@}��`6zu'2�F�Ȣ\�������-��X�N���DtK�_���D�X���\Zud�ͪ�1X,Xzb�k�o:���ll�l�wZ�S �ǽ;	M�?�$wg39vAn�,���rWôkB�3��>�5"���vK��s=���|ǒ{�p��r�pQ�s��;JI�X³�WLF�kz����n�w`9�E�"��o���^���T�ծY���mevʮ��ze菅|�ߵ,�@+e�f��ܟp㍮#��O�c�A�#�v����c+��t��b^1�e����2�@b'5�E6'�G*�'ć��9���Fii�/���>��gD]�lQI6���d�x|g�(BB�Q�׹�JP5&����jlv`�����N�Н?z7���'�`�J�z�d�s�	���Y����ʾ�g,7�^�b����ף��rk{��	�:ek[^b� X=}K�&I\,;�&�!,�)��\�l`��O��K��ٺ%�H��Oſ;�m���gP���67�'�9�US�F���5ŋ�M�m�ebbF����γ����RӾxd��ub�C	��T͏ఄ5�wq�6XbL��e���F=��&�N����I���#lE�J�洬��g��xM-Gr
%�h]��k)tM���c3��ԕ%N�5ޡ$�ߎ8;	\�)G2K�A�Ȟ-��;w����c#� 	���Y�ǫޗΆ��o%�<�yثydA����Ĺ�޿��0?qӗ>#�ƾ�g~v�A��Q[z�q{�|oGU
{E�b	���<����_��Ze|�R�L�p7��*����\�΂&����Y%��@Wдj�B{��+����1�~�.˪ ��!^/�^��f�<�	����	q���n��~Y5�����d�k��2��X������Nr���ọ؆�����e�����Ŷ�1�L�,ZT��y���[�}�}��jMu~{>�;��Ɇ��*ՠ��9!ք�L�S�p4	�+$Z�!����¨iv9�7�nu��KC�����0X��h�1�_18nĦ��[���@J)v$B����r��-=�/@��c�h���b]��=���+ϳ��RK���>�0����;&6��P��{'����aOTZ�6Td2�����a�v�I�j��K�:��#(��Ld��4��5 �G�!���zv �]�S+�p%�&uV�yZ��6`��,�٢ϘRnBѴ���F;�!H�SuY��',�6�ϯ�i�A�`j���efH�_�؏l ��dn� ���׀L�b�A���\��?�J4&�w9?��J�$��� } �N�3�e���[z�e͝�a1�G�+��܆KE�U�GA���#ڍ�Wa��#��q��-=�v�xʓ
.�O����Ml\=�M@���1
��]�:���ِ�@"4 6����QJ�+��Q#�t�S���MO%r����ZrH�V�vt�|�EF��*9f�x ڧ� 0#���(�/��~u��]
f,g?<%Q{��`򵀆v������:�f�Y�r���7�������L�z!G��4�o��C�4��W�� ����y�?Z�>��I;�N�B���*�3���h������u���/ɦ�}>��{d�/����y܎¨�a(�!��ߤ2�;�%��YP��T����u݇dMڌ����@?oOLR����#R4��JW��S0�3	�T�IA�r�$���`��X����o
�T?�u!r�Ɨ
h_Ec�ا+~6\yqgmԐqַ����)xp��K�
'Q�&�=O�M+��I0�2y
�%�/�Tb���L����O��0��r5`�GO7�C��|ۨ������3@gNl s>Ub�)�œѥ�Yyu"@y�0 �����9#1�R��4�P���c���8Yv����2��U��OάN;֞D��ME�,M��烶�W[H`e7������dM.O���)�^�+kq��O��Zna���K8����q�%B���� �4�X�F�7�C�˿7��6j��c��E!�v���|���B}F�QsN卼�a�~_?;�����X�TCn�`C�5U��3�mE������R�4��r�Y#�~���T��4fVYbE�7	w9Fyd�$͑�W(|�L�j�9W�j		�~��o�L�^�k�������d�Q��:�:��ƾ@n�z�_*�jؙ�y\7<��t�(������:?ߐ�p���&���R�ȗ�;�V��� ��)��+ee�S��Bt�����60�ii��ZZ����V�_U[�E�qԥ:nA��T�O���l��1�W�N2[�L��p�ԟSz,:��Hu1(�P�f����xmެwR��W�Ⴋ�Ypmvh���&µ��{��
��aD7�.'J����5w��EGa�&�#tS���f���5w|h�'g��b{"Q����/�jU�䂓�$�7�q��#��L�e�͏l�v�O¥�N�qz&��α!���$�:��h
��X���!*G��;��[�4�뱫~Q�+4�a����S�۔,��j4��f_�鸕EW���VD��d�.�Z�d>i/���f-�$}�fX�d��)�3آQ�b��Z��\W���[QD�L'e�Q��P�FIqY-���s T}����*�1���ra��(;X�E�+��`�۫�k���%�(Y)4a؝���(~y��C4:����(�>�(=8렾1:%"�@�[��U�%�i�U(Z㇧�z�de8�Bs�qf"'�31��l���=��EV����6�w��'�˹�C�� s�"�W!�3<���Yک�G!�*Q�W�1��	3�����mN�&�`l���ݳ��Եg˳�..��������Y���UpMNߧ46J���R!3J_9���/��:]��O$��*>?�1�������!�D&��C1Y�Uwպ\z7�"�������8c͒�f� �8��T�y�n�4F��r��f�߂`�?��~�bħ��4 򣦨��0Q9e�i.LHx���)Ku�h���V�
��IRe��%^��ޮ@�A�r�����E8	�>��u���,5�堽BK�h����n�L�ca-����tݒ��cv��S��S?H<����MpQ�HW�"���'HW�a�XMj����Gf�}^�;�|��v�ꇜ��ʿ���TG�I���.Y`�xeÞ	�,�M�-��_��_�џr>A��S)8(��ؖcw�,Mb�t�~�F�|O����tJT�e2/�Ǟr)����y�����e�!~�k~&���)��zM��m)�G��?��Z���xU��g^�&#!õf�#����r����J�!>�_~Ǭ�M��^9����3�6�ZG��R�3F�V�Ӳ�?{~�+3���z�����i��eI�.!�+�,��F) 	�1�������O��x�UX����aB�N`����B�_����ʼ~�X0E��NҀ�����0qބJ�]��������=�c�9�ʘw�Nd��̦��h¡E���d0{Z���3uI��զ~S��T6p�Aaj2g��c	�[�T{*<ӸՎ�?�}¼��B$��7�K�������:���]*�'��ʌtKa��ƿ����D���:c/Yw��j}�:���x�b�\$K"¼NM��]sȶ/�j�Q�|��� ��s��%,��3�ЦD}������B��g�@�����Ϝ2�$��S�_�f�d��]��}��>0lhݭ��^'P�ʹ_'Gдc �e0��U��VV�\S�S����Y�\L�O��=3H撁�ވ��P~�k�K��+�&es�l X0�Ŷ����H5$bU�(�kY7ih�^'+��u�Ɋ('��^Ƚ�2��!���q�e��|�'ڥ=�����*���Γ�g����ߡ��F���B욨?!iw����0�;+�ʼ�53s1�>�������޼�5p�d'�<�l/+�
_lי-7%p��8�, ��Cp@-����~��<P�n�AҼ~,)ᙼ�lD6�Y�)��i����0�=�!dt����eh�(�㎹=V0�k��U��gYcsnv��j�ǥ���o�B��M���Z�t_T�$��Tl $b�֊t��5��z۳��(��b:^�H�O���hG���'p��w�9�:{ec쑒��U�����d��W�{Y⑖��ӂȑN	d��<�OI��E������T���FY��׍o�I�Z��+��RQZ��J�qLo�����Os���QϢ���:���&_���#�!�����J�8�-��]�.v�BN��t�@����"g'@;��Q�a�i�)L���L�1�u�0@ǌ�y���ٱs`L��w7weH`�gxF�k�pSCč�_S�NP�O6;c����S���(j1bNN�)A_s�9ɍ�g^"I5�\��=@I<ũ ��^�HO���7�N��}1l���� �@��q����I�!��Bj�}߮+� �.p��4��\+ �ڮ���1oIţ0)H��1���jL���f���c��F�;�Ȱ��קO��1�)]k���6-P�|�NQ]��yB7 �(|���t4w%�V��j �-�-�s��"��MO͸��<�������K�f��� �'�!ɓ+��S3y�jğ�<�y�1�{���=�����qr�����K��K��4�]�� �����'�@6OMJ�!�M���vi~�8Y	6���@`�]��^Έ��)S�֮j �5�K[9�-�K���C�1�?䘬0�5oo��/�dW�o~�90N�^��ūon�"'�>u�?:�2O�)�. �ݘ�\YDsu-�o�-)�1°x��)�E���OJJ���nL龀��QoǠam�7l���xmPo�~P�����c��^�����q�.T:N&3��>-�
���a.�;��)i}�%����[�t V`#,��G�/Ǽ.���{3F�AͲ��^�3��O��)�h�6}X	���7���b�{�D^���+�~*��t�9�8	up\ۣcu�� �E�sˡ[8��MX�Ab[�1|U�þA��Hk֬��R9@��ʍ�V��-�(�-���V|�^`�p$�d-��&9 �M��?7�ޞ2ƛ�)�l���}��+��t�"?	m�v=�q���9��-Em�\ܢ*1�u������-\ʲ; ��fb�4Qm=�){͠�w��(��_�v׶�{�$��榘ob�Z��VZ%� ��=C8�]��BQ�L��->e�N�=�I�E|tN�h�f��^��mD�w� t\���i�_���gm�~�*���p=1�[�k�mP�;��|��)��om26eb���G�8�Nk�	O@L��?~�*U��}X��^=���NlhYdͷ��l����������Yc��sTo���"@��
��	��cK"kt1Ǆ4c]}�mڂ�&��ځt{�����Y�(e���/�f��Q�j������u���t�m�9v�vۍ�u�m4��9�*<'d��%�X������I�~��-9Н�̳?{mi��������u�g��x�w���`4"KB�WA�_y`��O5��>�?�eT�0q������ky�Y�ſL<+s�}x+���o�IE�`<�j;�@�""�쎝�� /q�$��,1�7Ɇǿ&�n�߇�H�K��Q���5f��l1���G�ly�J�	���+�9���D=[���ti�
���X����?�]�[�T3ѿ��y@ ��)���t�Ⴛ���tl�%b�i!����%��d![��$��gM�ϟN�Q2�ꏾ�16�<{LYB�n�U��ҕ	����� ֔�i��J�7?���L^&��n��
C�Za���*����&0�?j�A!���G	�n��C�vV�����'D���eV���b�)�����Zk�>��:߹� =%*<x��M�5�㐑�pvk�,@��qV�![����� ��5��%@8�K�(��
�@-��dY�V�CP���c�~z,�]�Y��d)=�k�<"9F��x��e�WimTH�3�0'�P �m�T��4
Q�L��2���>�T���ѤP?p�,�s�p2��(�c��_�MpƁ��[�;感�\˝�$c��) ��@�uns�$�������^��q� {)�a�<E�Q�U���z���k�6�?�r
N�#/'��\�<Ç�D��wl���3��K�x|�ǔ����C)�-�j8`�c�B	�Yk��4L��3�9��)�w�4�ڢc�H�n�Hs7-.կ C-��О��	�½x�W*d(v�̐b}8%��pށs��=ƴ�#ms�z�Ȱa�7cX|��%b���8)n+J� n��'F
�V3�/&���8
���b������@Y��s�3J��GIAz����/�n����ۀȰ൩�N�����AX�5���}-�hVM��z��Id�$�
n�׳G�T0��9R�b�䠂�M��)�\�[N�@����߈u��M��>���`%� t�Hݘ[����A���w���u��Q�CS����aM5���P�/"昸:`�ϕ%dvO �%�ۂ��b�<˔�],�[!��By;�b�%=�0�����������R�����Ɍ9�7����Lg�@(�y��͉��	��{�P���}
Zv��6��MR�6�f���~!eNa��ۏ��U�� m��@x��%ղKa�K}S���JM�`���A}h2�J���l�f��:��j�@���~��)�ovQ�\}}�[�vR�Y}�:�o?w#*!I(�o/V�^�o��V�Z���	���.��J�|��K;���� �SWSh�dKo����+$��Rv7,�l�|Z�ꎯC{�;��t͈r��x���s���MO&�4�I��_��f9�ϒ�#/��6@��U e���w�Q#�F�E����B�l�R�Ѭ"r�D�ͯ�:�4?�b���L�sV����y���N��]��
��%�Aff�r`j�S}�[����S	%�e@����F<rn�o�2��"���1�9L:C#l��4^]�=�Î:5����&|\���|3����	�Wv"��bc?T����q8����/��"����i��
��R���t'F�T�8�O�Dc����X_��*F��LS���&���¸n!��<1%����u�Wk�΢q��sfٰ��G-h=MAޚyl�9ZE��p}��˻��O!���t��y��#��r�kD���b'Q�aΥ�m·��>fK��"��9�x�'�Y��"|�g�a��䗳���,`6[�7��g�{���D�ţ��a��'��y�์}�_u��sw�ٱǯ]d��ѨG�=���`��I"�b*�f�Y�+�>R�:኿`>���F�1G�bMA5+_�KArhV�+������&�K�8뵘&o�g�m�X��};�����v�AjrU5��!	�TV� �������iw��%��LȬ����ij�Ɔ���:�k��I-Ց;��ךc_i�\a$�P5�
�ww4f|
w��
k�rÏ���N�燡��^)��������칷�� m�� ɵc`pP����4�Gv�'P^�Ĺ`FS_�*,5�w\�8%Wk��;�����-��};Y��<�'��lG9��|�Q�����ձ�>m�X�a�؃ �I�xɤ���N/)�[���VtJ���8��St�}�4[FQ+��G;����O@gxe���y��X�l{(�I8ܐ���]�׉7>f�~u�.p���*M0U�3�ű�uq�i�7��~fR"� �'e\��c,Ǉ`Q�HV���� �J����>�5F��8�m~��`��4ג<!��	��� �Z{��z��I�h�u:?����Ԁ{"�,�|��	��T}�/�����|!���;���}�<v�����*5�⁽'șrZWN�n
��S}sd~@���Rc�Jx�{�;��
�8׫�h;ޤ��b9�ѫX꒴�m�<K�}JY�	{q�]o.�M_���d����|M+$;���_қ4��h�T���E5g��X�^)C�,�O�v	������9Ⱦdb��@���:�iu��Ȱ����k�ڃuhT,�_|ڙ�F���pH�Ԯ/�"L�(rH�(\� �ڮǷF���<��Q��M�7/9 C}�;H#�ʀ �ϓ���EE��<CʨZ��L��#����:��7�Rj[�����l#���}]�p$s�XH�#&wU��Xx����d�_���(����\o]�� Z,*�0�ͦ+�� ����{ю���P^���������%f@9�>#�T���p��-f�������m��\�ۊ������%��p��q8�������Y[o��K�>cfԫ�{�^�c��q	ĉ��%���%�{ �Kx2����s�ǆ9�̤�+�:췡��n�Zi'��'F낮�_�Kz�"���~6��Ǌ�[�O��&���e:$�+mhI%����9��8L W\t?	��ui2�N��`�;l��E��"���N ������Û�g�d�V4.'�8;��Z��_��0%��?����oN��`��H��{=۩v����Gu��ص�0����ܾb��o�E\!�H{����f~5_������R?0�O�� �)���(�8[TI���1�rl����{�P�E5�Gږ��Ͽ7�6�;\*2F�����]ΧnǲZ�������Gї7��Y���=�<W���)��-pSnF5��i���"��噡�h�T�,�Yw�?�g�I�h6�w1����sˍf�{�#bN�RS��p~��R���8��Z'�M����@��<�{qr]iQ��I���ɥ�n�;䎴)��A��]]���Λ�X\699�3V�8��>�ەC3\��q�1S�l�־�5�tpo�$3ֶ��w^�����l�����.���S#���]�) ���e��cz�UQh���2�F�0�c~w�U���} �|O�gb��ʸ�b��e$_�`�6-��_m����N�k�q\�>�C����A�R9��bFv�ɞ�����쐓�	2�Q�>����&�`�Pu~��p�E����E�U`N����zKh�KIP۰b��db�θ��AW.v�u�QGt3����^ҁ��q���� ��1��Fٰ��n./,띜�O6���5���!P���vK:�/���dfbt�Y����� ���C=�m8��_pZ��<��2br�Y������2"3BƗ�+���Mm�:�j����K�C�����ZW�����G:�����RRo���Ƶ�j5툚W�R�����WxI�����C�R��-՟��aH��F��h�j:���2��z�?�Mu�����T�N��
O�ZYʿ=�Ds~���|�}F\�ìxOY����=l�������\�!L���5,�{B���7Ƅ6�Q�uS��t�߼7�i'�;��|��;LX`m=_9�c�?aX���o:���=�g�I��N5?+��W����SH!.T�k��ۘ*�X���ʃ�KU��M�ɉ�Ѣ�#*���q�x=�g �^�J�0�M: F�|ꉦ�.���yg�t}�����2�� �F���/WI�g �x=����<�g��X� +��=p�>� �|������������,��c���	I��o+`��b��?a�D�J�D�HOݴ�?�q�H�a;`gg�����u������?�#L��Ëk�
e�i�=�-�����M�΃����)�:�cNnZ�%�J�9��?�U�2�zXD<k	cq7�!�&��&��{|��S3?�y)bس��c��+�ˀ˲���$<�7
{+k���o�@��7��*��&�Ʈ��˶>���BĐĹ�@���$3/�?��D�jH�+tQ�/���1(�r��h�Q����J�)O<��s��*�@8DWm:�8�[O)_я�zdc��[k3�e}��_:�R<ܗ4�g�}>�͗�.~�t� ���"�r�FKHD�*=�NSp�GhQۃPr���9��Y)��-�갳@-Q1�=�O�`�/��9m*�	�J���I�1x�����R�Z����rA��H|��`{a'Es�!��E׏��B(q 11x�j h��BC#��l`�.���%�O%I��L q�wJ�B�k��g~��2��(!ܚc���8��=���MX� o(l�R�����&���tv�[�w�6)����g�@����t�-���_���~���A�n(�ToGb����!�@��W���p����O}T�Hii�b����h��v\ʅ�4��J�����剝%x�K��EÖkkV1��O�j����>d�+�8�L��rN����&-I�mH6��~��������g_�La\����������3���CR���Rݾ���?VJ=�Nȹ�36,��o;^��b?l�^<�r��V�@���P<��1��YJ{�Hܒ菬9b�u^�t��+t~�#��G+;$�~��<T��d��Y=��~��i�ۊ�����a��+q����0:�+�񠬓�'z�7�) �ؑ��M���A�+c�t�ֻ�FS�f���-��D�#J(JҐ�4sS��1�Cap3� �8b�B�����������'�O�O	��`0z��r^�����rq��o���~D�:�j,$����y��,���Ϳ�>�J�h�&��;��|\�*��{�p񛫂�gz��[�U����W�F aJ�R*���2fV.&]ɣҊѕ���w�B��`)����B��=BaP9j�s�)�[�Vj
fJ:'���ڕ�;��/�[�ѱ��r��+,W�\���]�
�bF���CY�.��y��::��'1m��#ρ4�s��ng�)Qz8�_����za�d�]�� ˊ#�B���s-g�mM_2(5�|���Z���^ߑ��Kx�bRTR��#��:��M�6��r�t �I6] �!n���rSz��oj�Nʖ�#*�"E�W.VG%V����Ԃ����i�+��I���.���BG>�3U���Ic�
�}�Q��k>׋NݺG)21�h��3h<}�e�6\r ׻J���^�9��(�d6�֞��q^F�&���@�Y�)`��U�T�sY�:`�Ԓy��1���>-�'ȑq���"�u��ѽc�3v�]S�3�^��}���ƛ,�j��-jS��H�b����]��]� &I�2�ۧ/cs�_g��Ǣ�6<@��멣�y�0
 ��1�P�����P���m��G���3��s{k���X^i��]�,-��_��C�~�A{�ɩq��	�^d-L�yW�Tg�Gb������I�T�lTS��O|Rto��������=���Њ�u��tj�פ���v�Sr@�}8G�sÓT�� -S����"K��Z�ȣ0�\VU�-�.?8d��'P#�!�ׇ��kG��rT?�c%C��A�S��K��^����k��UJ(������jz�ϊ`n�X�6F��H�#���ؓ��Iؒ�5��6��Xv�r���<bL�"_�9���i�Za���Wq�`��i4��	&��G�K�b�-I��w�&�@����(K��z�?�ܵ�y���Jhnگl�rl��iK��4�y�$�r��$%p'�ڧ�f�W��akρ�M�Ht�3�ᔙ!P�5�8|������~�
2�f�\�*�pE'��43�m���v��S���8 �+�N�f�]ã!���S�A�C.c� ���^>�}JaPӧ�b�]j���AT�-,R����:�V��:�<� ��ΰ^ud�G��v���4�2���,�l�|�)�*�F-=�E��Pq0�Btnd���U�e��b�J�;��	tjC�)Ä�c��5n��z�T`��g������A#A� Jn��ՀS�[��ι����1��&YO�!�{�ʣ#�T�r!���w`�`\93�>�rJ\����u���(d@�n\�؊�67���^A�[�p �P��	!�.�GQ~""����%v0CF�ӑEbۍ�X�:���oh.��0����>�����d�ǜ:���WI���g?_i��yW��a�)�-CF��Nǂ[x��A�>�IeR&����2U��z������έr�E���͈Pz�W��7 Z�32����T�u��|����݁	�(�z�Z6��\rr�#R���[�+y���u>����w�Q)�L9�o��[,.��t��Җ�s~l'3qF�'I	�{�aiE�A�j#E�|�h�. M�rF�n����?β{j�yo4t=���O�؆�d�T>M�忛�iq'�f���p\]C�`2&,�ߍ���'i��E�$��_b͌��sZ.�]qpF�����~1�C�S�%����j�=�YB %zɡF2�a���θ|��C�x�wa���ӫ (�x�L��jl̲�*���c؜w�!vGyj�-fT{�R��;İ�������]2�F��M�4 �Ӭ�$��Ja�������Y��<Y�o��c-0P�:q����o��y^n����Sښ!C��%��ρ��=7G[I۹V��wV�+��|�Oh�H�ip�(�G��՛�������s0�$�*.F˯��%]2���,A&�W;��� l�4��o�;��w��eڋ��!	/C���uE�S{�"`ѡ����	_1����~��	?�i��'�
�~+.Ot�ٿwj��.oa�idf�̥:���I0��2����0�2��7������[�/��zz�P+W�f��wp��1Wm����o���a ���Mf4�H���,�?�X�i�:����Z�'0"K�r�80K(2�C�&�N[^��Ex�5).E��yA��|����P�8� Bi��>����x��q�B���$0X=�"���k�|�*������+ʋӱ�4�|g���ד-9;����n̸e��mm�$������~0�����e��_��Ϟ��#����&wg^ǲ�P���i��~���T�<�)&=����t5#cH,dk�#�H��v���5s.N���qo�~����j�n�^$�oc��%	UӸ��Q�,��5E���M�W��r���%fF��X�MzX)���="���Ad_������N	���-rwT\���At{/�ҿ�zE���;*n������zXc�0x�l���r��U:�ܩ@n ���!��xnrNB���;Q� ��i���)��Ӣz�Zӈ���-j����*�%�ꗩ�0�=]�:�s�%��FR�`/���Fo�f4�_z�٭��k)���8wwI�A���T�����vkb�]��9m�UR�����-HSH��F��H�h�=gV����8����yNo�@Ӳ�M����n�тR0O�3���_���2�ˀ�ѴKS�O���ٺ1Ւ�����+Φ9`#�)������:6H៯x^�_�ok�[�9�o�s:#?�y�����8�Zw��"�˱�ԯ�qr��B�Q�gV��뿉L��G��=��R�hϛL �,��Y�QE`��A]�v[��s=ɷo��OU��r�0{l���BI.0rz5�҄�O�=��z�DH������{�������Ϥ�ֈ��k3���FYc�4-B�b/no!�v�℞و�3+�1��GZ�޶����*�V�n�K�P���5�J�sp��1�Jy�CR��,m�<�F�Ɇ�ي�O�{}�Y����.�Z�1�*շq܌�X}ϥ�y�T�t�a)�t�M>����εB����\t"o�q1K���r�o���>7g7���[��	��^���	b�>�T��n��J3�|�c#!V��OG`��(���e�dH��7��p�K֞��'D���6(�ފ�ݞ6�8�0�nT(�2އ?�ᚯ��-��������H�-Ėd�ģ�>|nQt	IX@����M�R�E�ڔ/H�Ѣ��^W؂rz"VC�t�U{�vJ� �G���&�� S ��^����%��`<�Ik���T���H?�́�@�ĕH��ڇb����l���H8������ލc���"(���La=̲����Ec|���ډ����B���9j����(���Xw��t��0�
��Y�|���0���F�Ñ�kT�C���H{�;F�l�\q�p�\�|P?Dg��Ə�~���>i<�3׈l�@�K� �K��I�Qhn��=d�+��j# ~��l{�R��C����m��/��g���Y��yaS�0?�5�1�q�*LZN�f	C�S1��
M��~�%W�}t����]��7�"��R�~�+~�&�
�ҵå�)/��B����ҵy�8���}��D/v�Ccg�\�Z� �J�9���:�*�1����<���{�-���4�s�,D�n�g�!��
�)^��g��ي��'��R-�ώw�#�O�"���B�hI5~ ���Γ,X�b�Hר(oC���\�.�L���s;EsM�V��`�p��d3I�'νA�O��<S=]�=��IW�Y��o_%���G��d�tf�
�+��Y�mMO�P)Jg�.F($;���֞�Ihl��:38����)?��E)��<v���x�u�Q,:q�"7M�Do4.���0>��(8[���.=��]}}bٓٵ*����$��������]Kz����VwZ?&fG��$ޱ����s�����j؁)[[2�6���9f�~�QA�s���6{w�w��>u�5AH� ��5��6��m�h����B���D�M�ٍAʤk�s�N��!f��3���	��a1�8$�5.�Vq���uU�N�vV�L�-t��mL��q!�*jz8(�!�Ե�(�Vl��!�I��o�`#'��A�y������0�d��{��QO ֜]є� =��L@���#p��<��B�Rr��1o��Y��L�C�]'�yV][�Y�l��b�
/��ΕL�IG8!�)�QΏ��������O���ȳ��Y]����I~�S��r�dÎ(��b�o����ؿ�kbEA�Cv;i<#�p�����gqN!�CVH���G���̐v)����i�H۱`�g1�8�N����k�p���V>xGamH���KG��Z|n�a�	-ɰe3���w��T�O��,�}�+Hv���4�������NT4H�2��e�U�@�zj,�,2��d~�vi qC��݆�i�-R�'˭�q�pJ�	w)	���{'���,�s �	>$��w�8�#zI�r�sG�Ҁ ˨�躨�!�E�g�)Q�?��^Zb�ҝ�6�vgG���Ow|�E2l@�­���݉�7�ŉ�]���+�g�lb鬶V`���/K�>�`�#�} C�ε�����Q��H�O�cؿn�D��@H� ��e[G�	P�|)\V��}g�h��"���HÁ�L���q/�����]6�
}	,����a1m�����u
1.�۩�Ey]i<8"�@x��� �vC#<��*/�v�k�-H 8n�'�	�4]�_�hH�%/�W=�O��ZkTZ�|ވ'@������[�L�|Qp���#��&$T*ƈ駒��%���ȃ�EX�:w� !x�!�WlSq�J�FY�D�DS�w�';wk0�����='����grFY^U���P��g�r"�����L��nK��Pe��oʍ~s�S��r�.}5IB�OI����ϖ��AZ#��ϵ3ǉU[�����>A?;�u?�I�i�{~�mi�G!&'�����
|��i+Vg^:KN
��:һ�Vpl)����b�V��hW����.up�J��l����x�[nO̀+61&�*�v'\�����)�+��R&�n�8�hf�,E��]6�R5�{��Q�i�Պ���,�Hʺ@fa���2�
�!�|nj\a���v&'��|rE3��s͝Mf��`Iʌ���nr�ʃ�$�P�	u�Z[XJ�@��Ѩ��d㼕�3v�C/m�8l 2�M���C>T%c$�:���ΓT�E���m�K�p��Ԭ�G'��%���g��D	�9#�3�x�Fv�=i��@�b��)�L+��*1c�n�v
��׿����p4L����|��-ao֞�ZZ�]���\>;�y�+��1 ǂ�(���/pc��Z��Sv����M�h�X)a)HB��A�jQ�X�)��ԕ����w�k��z�+Q!��fif?��k�cfk�@ �~�Cw7���hy�����@�����"[�b�\�C"�����%���c�-��9R+o!���Q�vF��L�Ź��4}i��Ǽ潌�����A��d�^�#���x&��%G4��Q��j�7.�ϗ�B�j'C��2]�JSa��Nf�4�����ƣ�G�z�xg�FZ*>k���ƪ�9
�H�:�`�\O�^���lK&2�Z����-��Pr���f*r!�X�y���2B�xq>��?5��x}�5���l7����v�Ud�!�����%���RK���ƽ�b��P�Μ��N�)�Ʌ�ˏTˆ�oE���/<C%����t�JjEɉ�^~�}2%�z �}3�a>�c$?�!���ye'�$����[4�*8��ly��L`.��8��P�֧��/��}���ھ��#!������*�A��K����b �ٗ3}�R!>,��~:�����㷨��5G�e�%�c+�{��U���ڗ�82�]j��;�ͺV}���x��~�%�Mmm�W�x\��'?�*i���?�von��
�ϰ@y��@���/��2;-.�j�n���)�#�#��K��W�u�B��SqF��9+��8�S.D&���T���v���H�RZú
�2��V��[	s-t�4j_�0�̖%=\5�{�[%2*B�̆V������DC��3s�:I	g�S�
����W��*`��ð�baL�F	
I!��_>��d��0�,��È��6ė5v|�7�W��N�dA*b��4�V#q~�+r�hc_E�H�;�P��U��l/Tqڽ�P[g|�@��o�GX{*؆��SK����T������*�M�t8H�L�����P��)��$����8N���Ɉ�[���t��#k	��v���-�u�ƻô��,���Yx�Jm�`�z��ms�6�𬥈VOS\�/*�w�%G�9�<�au�6L@�=�����=9lD?�{M�c��V3* p� !����ޖN�A�@8��'T��%�)�1a7tj73>��"7<��H���o��Ӌ��gj+~	��[��L�ґӚ�iK�tk�9�Nj��U	7�+w/6���w�7��~��K�¢7��-�D��f��e�Λ.z����n
����>gP�,�3��O!gz�*[��l��� +��'��`�Wj6�����>�.��f3;�o�n0l��XuFe❮I�k��xT���H�Wp!6Is���vL�'���nw,.����ɲ�Bŧk�IQܘ�����S�3���Ob��@Oф��z�vZ�` �QY´���6J�+
ѿ����� ��]X	��a\�7j�+�Y��-�⼑H�m��[�'}����H� ��`���k����(&eq�*��7��\��/��R,$K�1��)Ж����|ؚ�[pU��A�{x�!���*��.�'9�_5q��V�dT)�G�k�]�vA��'*F6;���$��Dš�dHy����q��j�����5:MZ���()<V���c���q�����{_���rU1���Y�?Wa�[j]S<�츇,+J�,�ڌ�,%��6%)ĳ�ͨ��Ic,�����y�����Qՠy�u�f�S�׀X1�j4ljn��g8��\�ޢ%RڒX�̗ 2���om���Wm���>v�����,m)aP(]� �I���l�Ī��*!�_l��%�����,'�Wf��'��(�_E�t1�9�e�n��YJ���bko��
��m렭�h����c���5Jqm@V��ΰet�I��@M����Dן)Covݪn\�,8��6�i�cK�Nsb ��|2��ȭ�A<i�i�4h�2\l��G-���y�cŎ	��0'�����]���?�t���1��y7Y,�u�h[d�~P�����ki8�0�\4��s3��V��p�-� �CK���-^o\��fɭ���L+\9+A(���2���A��>�%.P;ºԉ�3�A�XN�o����-�%Q8�6�'N0C�+㤮����d�{`,��h_�?z�6G��0ɀVԭU_���U��ci�`��9N�׶�*�~���z艕L_����9+h@I�����g��vaQ�0���m�a`��MN�Nu�y��rw�@;o�Z����_����L䶥}��>�OˬA��`��R��~�"���&b��&j���m������#q�]���g
�>�������YB5~]�͞�%ޭq6\ZqW*`Dq����IY�&O	�|ON)�j{1g�?�
�tvgb��as����z�[F�����
Jl9�20�N�����[������|ݟ �P<�,1,,�*@���
� �2��bRՒ�:�O��еeZ��ˎ����SZ��a�s9�]ʏ��hH�D>�#�Xm7��1�����pK:��^8X�d�G�]|^����ss���
���z���n���l��3veM�����B�aq1���X�A�z�����^?j�O1�nB5䰋�;�Q�*���)��B0P^_ߝ'B��yVQ����`���Ɣ�$�P�!���_}��Wu��F���}v־��#���uAQM��.�݆7����7X�&�^�RE��x����rti�L��7m�\1�����������޴�&%�͂�����B�y����,��=�VW��G�NHK��L}�J��M��t{���+�i׃�J��Lv�X
ޘ������;�^%:@Fj18��L��E�|�uGS�
h��NiM|L�=u.hh�ć>A�����E�!���!^����n��9	{���pYЀ($����	I��X�V��k�(�m�{>6�
�A_�8�o��&�=����_���g��M7@���3��;\L�AU�R��fȺ��=�����"u�<�S>���p������2+�/�t�=�˽ڂ�Č��>M��?��Tߣ"<��ʪh�/֐�p}R��u}�Zeг.�"8��-�ӥ���avRL<�Kya#�A(I`�~ԝ0pULI�S���b(�����rk��H����]�TA�B;y�,ؾ��';�.C��x���&,��ރ����_�U�?�]�Է���p_-��ZJ������N�m�m�d�9SU�f���0Y���E �lGv�Ŀ_8���L�۫���PqG�"1�����7�s�%}��=)���9���xiT�i r���v�3"CCTqDX�E�DF�Ko<�,3��\2��諢Db�e\1����<� �'�@]�1�^ץ	��0@f�>�o�G��0��@���8��[?)�LYL���r���T_��6ƌ�J���h�b��(`Uj���OW����z�q�#h�!�����-O�ܫ��6d�ϟt��R�2J�0��eNE���i�B���g,	���������É�ul����U6���UGcjG�G��I0e0�-�������6B���7S�@CP_�$/{W%U���=ŪQ��3����[��K<�g6N$�Rp�
��t� +�L�5�K�H�Ko�`���H��eF��"��YB�ՠ���K1�S�i�Y <�"�~k��ì摾�l�igT%3���S*�������򻇬L�8H��B�D���D��b���y�:+S�#ҭN�
�b��z�ٞBI�$��G��/ތ0ǉ->S�\>I	�jƣ��rѫ�[���� ��IR݂`I�cfE��H���eޞ��!wc�$��C�/8��#R�w,�K,��8�H��c[*/����U��	�I��sG�2���	.���&��4Y�|v]�9��[)|i_� Z�;�`?��v^�JƗonB���S�)C���Զ��܄?[D_W��@P�V��ű�aP}�߬�c�a��-#ZRm�ևpo�z��pP�E� �c�\�k|%ؔ��'�֞wj�Yi<����{�[&�q��f���Τ2�#ʴ5u"�ʰ�l�W]�0ʠόd�E>x�j�#j��Ɯ=�8*�����]���<�@��_��N��HQS��^�s��*�~t�JK�8�t�Q-(/�-)���QI����髉w<�9=��Ma;J.�<�[��0�����,V%ϊ����`���P�O�#J�/"QyBt|���N:?�7U�p����G�vA���x�&6�M���]����˘$A��A��A���&2pZ�aͣLm�q/�)Bl�"��ufSm�/%��g�,6��]��*�����N���l�<8�q_��3eD,�O�?��6���p�[�ꬍ��S4�1���k}�Z��;�2c4n���Qm����h~-=	�58��h���*��]z>��ʕ�VL���W�[.��v��>`p��[iNQe?����Gb�g��ի��4e��X�ir�U��A��U0�;���~6�b�q�s�d�63=��;��^�{�h�6As}��}`����2��l��=#De��<{q� �MGt�}��(�Y��t��1�)����s������g��� ��=��kI�m�MӀ������!�$�w��	�1I�,�g�NYʨ/�T�8���h-�aX�`�ɚ�l� �e�%
�V"Q� �2te�qHM݇O<v����fa�r���}P��}*�o ����o��&Ѳ��IE�����*���߷�͂)Bn�H�����z�!̲S���h�h/^����"֒�D4�D~ʩ�J[;د�tW��'��_%��7�K}��m"k^�|-u��dS��������,.�Oé'���gG��]��a/��~쯶:b���X����젗�B�=Na!���p���Z������ɧ��-�#��؍�t&�
[�l�l��>jo��Ƃ��RN�Ri��ri������S�!+��^HIhjy�h�R�ii.�>�XbDt�X�Ľ�:I�W�̴��E1�vPp)g(kw�.v����D)+���9X�e!��X*9����*Em8LT��% ��{���Ӳ����M5oW�8����Y�l���KZ��Aa�|�rIp��H��}�L(;xg3_UIϯh�r|��S?�	�є���A�?Z����a�-�k\���E�8u�D���N�H]r��R�aLZ����
��[�4g��'�T�s�z��$��Kp\y��uk��mo��nv�����$�و7gM��ͭW;}i%���>�bν�҉�x������?��>S�Do�vD�mGz;,ƴ��c�g��FHa���-P���M�ό�"HD���t-�B�!�� �#���ׯ;��gظ��aS��Y=��kaÏ��~��*%�h���`ĚC�5����#6d#,%��%�L-���7a�#j�кU����ǉ�"��a� yV�Ec�q�t�	.^���H]�*+T��Qo}ۨ��X�Ak#^��K��cm9F9�_S����H�h���F��Rj�
ܦK�h̕��[섚�z�2� �y`X7��b|l����Հ������|l��" �!�g�6��;2nª�u��,�W���&�'��M�w��j(k�|c����#vA.4l�g�<d7�А}%���~A�$���^���&��M?��ӷ�4��t�_�!���ʡ�v��2T�C۽��/ŏ�琊�
����f9V��t�8e��}0���D��kk5�$~i��M�o�Pl\a���`%,'ޙQ������_��R�!���u� (�Ap���.(�����G�Y�͸�q��{
a@ߣ!�~﬍��tHQR�v��Y��_1�T�M�C'Q�ݛ�Y�{� 
�N~4�ƒ�W�$�q��a�����\���U�օN���q����`�Dg|?��Nn0)�"��CG�*hO��E�Ad�L_W_�M�,��v��G����>���Ս��.�Y\	���Q.8]���Z��ѻ�� ���*���	�b\��<2�p���͎;5D�$$�#:�/U�n�Ф�;_bU��e2?����s��z�L��+�ן�Q�'���e�
��^wY*�#��\l?�(L#_Q0(��	�ν'�=�g�Ĕ���q���J}_���x��
6��_�N��<��_)�\xw���*��}�PG!��^[���k�fh4�Y��U�ƅ�"�m+t<��ktB)��B��}4o{|��R۷Q[�V0H.�jYMy�O$w���"�@��ۇ:��.D���>�T�r#J4���c~K}�t�+�%B��۸Z�l4���abs��6ld�pVaFŬ,����w,� �v��E����NndF�7�����\'Ed����T�gqf�lZ����s�&��x��2��?�m��Z�p�	q��:�?�9���p��2+�E�:�E�����~D�^�A�f0\V�
e5��>��B���^%H����wܗ�<D���ǋr�.��g���H ����'�\��̰,����ps�hӾb/�M�KWL$��@}����ݑ'�_9Η�o��#�N�S�#=����qiUvȱq��"�8�k6�w<j�M�ز�X��I$�����䨉2%�C@l%Ԧ��m�Uw>�cF��8m꼩��d�w�u�DO�N��0�|���9���ƤG:����b�KXK�3���8��5GW��܈"}��y�Qv5e�9�Wd�4���c��{�ݲԎFb��ye橅�&�N�6�9�%B_`mf�E�Pa�nXܘG4����n@NJN;u���N����Q��~h'(�X�NW�=��g�� ^˺]�p��J@ܬ�M�^e����,T�1Ӑ�u��IK���j?�����ä���Ͼ;�_/.ʈ��CB�t��'C|'kc�qh7��}�emw�kS�RDO˳pv(�9�0�6�����-�yl-o�#�(������uK�2���J��{��,};�ٶL  ���! ԂT�K4��TH��|y�	�aq��l��C���0�#텄fgP{���vq���0��>߾�X�X�	1��y��ox���/g�>}㕎�DbzqA���b$��D���Ur��	n��j���:�lZ�o�v���M܆� ʲ��vO�%�3�R��B��f�\?3��Ga�M�)��D8�K8�$�	6���ܮ6U(�Nc��|K��/�ǯ;�+,1L���_�����$�ƿ�m����o�������UeT�妠�!����M%�h��0�ҹ�G��{O<F��I��O�"S~Ư�W*���~��@�>�-�w۩�<,n�<�v�z��8�)�gb�\3B6�ԙ㮐9�,JvѶ��f��.�_)kNd8I��=&�T�~e��+����q*�:�"Yʞe>"-������)H�w֥F��J�d!���������I�ZPv	vn�����F�;�5:e;���w�톚���m�KEC�g㚹y�D��%#�FE�6��o��j*�ߝn�梠>�*E]��"ٟ|��$�$�
��9%"��Q^�+=;?j�~ IR����?�a~p �ō���(>����ʭ+����68�z��\0�	��a�×wsY�b��=�9�l��|j�y��\)�H�j���f�_�-M�E,�E/pJ��S�.�9�fCߊ��T�FN��a��ܰ[�Iܤ�\Bq��F�&^���*ۻyh�*���'�Q]��ͧ7H�	�hJk�p�Ş��;���Hd���X'C����0e��#��G��˛��[ݝ��L505gК�;Qɽ�3T�g��A�����'���îB;D^�d�x8���6��EP���2�7:��f543B�#��*\�ժ���͆4��̴��F�8�L��
6��N;�#���G3.����Q)n0�P�+C&��)x�+3HA�J��®�sA[���Jv]�1m���tϝ�'����<�K�Uy�!<�����g��o��TWջśQ�)`��U�X\W�����ӾғCJr�nK��QD{}���Ɓ���}�LB[̩�\p�2a�u�"~h�J�3�"���ߨU#G]�-����aڟ�2S��fh.O��E�_e�¿|�k�k`���"S�:3{��
'H���y��N�#�	��ܡ�v�i� ol�&��p�m��F����m������� ��g�j ���8d��粫c����Y�^���Y���m�97�^�;HA;�{�P��偲e����_��������5�H�����HEz���4��F�Q���Q.���5!XOb�3�{D��K���a�����\�E�P�dLx#O�Gw|��=��2�o:����T�h����(ʣ��F볺��q����L��W���+T��MԈ���8��b�Y�w���x|�G�UŞ�U��n�7���z��R?(������5�MZ�����-���?mR���*AOu�8����d�)���h�;�y��-N9ڞ\�hG��d�s�#>�̪#�����5�ۉ^�.�G����H�=�&j�Nj�[3��u�|��R��
Vm�F��`h� Ǟ�,w��ܰ��1���D��^��
f�4nW��"��������9DY{(m{Q��S	p/��p����k�����5���_��ub8��Vă	���F?3Y)����v+��k ��V�������� �f�[_�)�� T�ן�Z68l�R)��ޙ�� ��]��@^v�����N��{^#��aQt��c�CIio������C'�IU+c�j��{#@�/�<��[���	#w�P����پ�Fగ�	��%`�ƺ
�>�u���&/K<�&����S-� ̠�����=���OI/V��J�,B(9:�nSw���pSIxՂ2��Yw�<�a�j�D�'�m�����+sӓ����+H2��U���ؚaK���
of���N�p���|���^��f��a���x�-�{4ܦCX�$c,$�+�U/T�n!ٿ�����h�9"��K%�w���<��a�G��4@��F���O�����;dh�����(�ӯ�q��*�1���׋�ﶒ^_«��������V^���uX�m~k0PT� }�1��u���}3��K�%}�1n*�qҶG�?�����)·���#մw�"/7�	�7�;3�]�E8)2ח�pet�`H+�����N��=rW������FN0I�M��M��50xy wd�m#q�	>R�I�b��J4�S�F��ɞ�q ��V�m|�l��o�Q�i("֭풾�3���͊��\��\��zP�y�[���ܧ	��8��Mt{��L���d��o�3�j>F�9쮮�c5W{XӀA����������27�ѷϹ�V9L�DN��2wN����h2R���l���ęUQ�Q��/����$0�2'��pK�8�a����967Pݮ�~� �.��{�^B��$G���e�b�;�����L��J��W�+�K�|� ��;~��b�ZT��C�.#*���6�4�,����\s@�qF̻	{ۮŇ�����!��zfL����V��7����j�gH�g�� ���c�ꖷc�lH��"C��.�S��q�)��28�ȩD�qᣄO�=����Z�y�ve�R���r�d/����ž�ǅ���z��o���A��ެK��Ě�{#F�tyyQ�ӗ�Q�(�< �!�"��wճu���F^k�^���-�Le�)=�7�dQ������4 7^2e9��wp�pI[�ު��Oj&�t�|#a�tix���V���c���=t�GY���4�k�\!y}3Ѻ
�J���6���#���8of�kcƋ�װ!��JFu&6�o� 4�f���5Y�nڭ�l�Y�AKSM��Z��(9�c����v)mb�8,<�a3R� ��eFn�b;�ɞ?�L�0i?����i�
�S�]7��?T�ȋ*���j�o��=�f8�_�����(��Ya�P��������#7�Y�ƕz]�S[M�b�]6�;�X�C����l���+��_� �����8ՏK2p�Vf?�zGC窢`�����Q#�5���L�е6J�<js�n��a�&SH�%�Yޚ���jj��>�b�.���6�b߯�n	b��,���]�sIǻt��{�g����1.I* Y'�0,x�wvԘrҽ�3ћ���I}k��챲ωV�/�����6Rq�|zcx�Zz�qܣ+�P�Kqy3?,� w6_�S����"T&@D��%���z�?�:;}�uo�x�mE]捊��"��g|ǚ��-����l�F�T_�m��]�Denu�I,j�9#�E��9�n\�?����;�֗#�1�B����6[��O��c�M�B+?�-�@�����Ǭ�'�{k�~N֎��ߏZ�i��ʪ�3$�~���X��#R��[���_��@�`�?i&�_z�ER�V�x�[8X�P�#��d���4 ����߿�'��]��OY]��{�a��;�V�Cc/�m��.�>7m�Eˮ�Υ�����H]�Y�R�_b��p=`�s����#�_�8����B�|�|T���nF�N*�tf���N������v/n%1l���YeM4��-�d:n'��gϪ�Oá
���}�[y��c�ඞ.D�#�T���7�&�7�剜|B�4�D������Bs�K�<�|�v=A�[�,����(�	�12Y��,K�a���GJ��\�ӂ�E������r��Ǫl礚�ز���aKߋ�����
!������:H@Il�;Z̅��'�݆8;z7�E''U��3����m��W��"׾6�=��/d��o�����AS"���I�Vq��Olve^~��º�������W\���[��os�6�{����<$���w��� ƨ�/m�Α��⿍Ȥ�]uzZ�6o�o��c���ߞ"�wקҥ��g�P�Jsf�@R�7�����q*��}o*�E����/��vĽR+��R�I�h�D=����#sϔ�pp'�DQ&�,T��D49֣̀�<��K]�H�f�l�P��2�zv~�']y��C&寓�ܽ�cwdğ����l��k�L.K����d&I4�r������:`/}�����H�ZS�c��1���4�|�0#�J�q��1,�d9����0z�K��/��z�򂌇W_��H����=����|����@#�ܬ�d&J�p�F�����/�ĸ�ގ)��>2f��i��%��C�\h��aB�7F�\-Ÿ���y�XtfRQ";غ���A[��-0ۨ��]G|ƔP�փ�u8����S�=A��O}�@�9w��[���0y��S��=E�׵4]�p涄���~�%π���i��ݣS�6��1Φ�$���
M2�Ɏ��I���j���5%��k�P�g��A@ih0x�����~R��N}:�^�����=���r��0�
�E�F�^����LM��}��FO�:�;v��Q�ĤgZFf�tz�9!^bGo4%�����|v��\��t����U��������}����&8��R��j9��Y𤋷o���]#<k��@�@E�䈌J�#߸��VZp^�PĘ���.,�re��f��j*L�joD��IM�jϔ�D����Lvi��rP��׊)�ۓ�,HI��sk��	؁��x�����0 f��#\
��Aq��0�f]fgޔAA��(�n$�{�O}����-�'zs���5����bS��K�$��ڴ�H�~֫��~��Oˤ��Q�#R��m��n�T*˦N�	6��<=�$c9��u<�u0lB��v�,�'�L��KQ�p��[�W����hjsSa�57�"�
�l� +�vkD,��k��[��~��c�x��z��Mw����#c2�Hp�O.T�-�#z#�=�˜@�8�в������5+�u�`N��N��(��m��A:Q�=�
ea\�ۀ�[�55��>e瀔C���>8������O^Rv�h�r��E:,2�����H
cz`�P�μ(!ʮ�6��ּ�{�wK�H�%q��GH��|��Y�����C���J�hآ�(�=� 1�*O�;��S�r�-S~�L���8��Q�Ĭ'�j��Juy Q�E�9s/ȇ	���h�)�*��y7��t��)�t��v���	K������>@���A;.!1$7
���q��� ׌8J��y_>�;�6{�w�b`ݲ��Ō7qMp�dآ�m����f6Z���-~6]k""�0� �4U"F���$�5�枫U����|���5�h�wŊ��6^F�jbcw�P���;m]Vr&�^jFŊ��#h��B� �H�J��'`UG��1��,�V��E?����M.4?m�[��дI��n��8�����MR&�Ł}+q��D���|7E�Bw��J� �Ʈ9Íy���>q@�M���:�=�Ė�S�
��˜% ��|O/��`��rjx�6,����s�7����>���f��^H��@��arq�=�'~e-���b_��0 ����Ir����� ���tU�]�Qџ�0=<�S������?s��[���*Q��
G��]t�%v�����p�z�� ��[x��]ڭt��pC>3;"������qrw���I��K�I����Z;��K��>U�b����9'���7r��h�{���O�)����ĥ��2y���mͻg�g������� ���SQق!��j(�G6vYh�]-���&i���pi��c7��K�=���}�S&��S�AI��V�.`^��~�Ԇrf��^I����&|/����b���·W�d�z{����0p�3�{]O��-u�{���b�y�eb�����K�'>^��WA�q��]�E���F7�����X�(sHBq�(,?�;�ZbQ������v�J_lj� }J��_��{P�-�,@��4�˱�X���kw����o����\i��<J�O�Sr�L7���ΏD@jй��8N�Ę����k__r�s�%���*�D���d�� g���@I,�o��N�׷M�Y�X��'�j�r�p���Gȫ]����MVH-�@���G�*���-��V����r��$r�Z��}�~����G�DȷBi���=CJg{��6�"��Y��vݕ�-�ӋQ �9�a	�%
�2��0��V�~NG�RQ��L.� Вԝ��1�!Υ��2u<�aˁ\�	�Vs���U��I�����]h[K���3Hj����28T)�]j�V�U.��5:bR�č���0�����@��Ȋ��QV	(ݩ[QH�Qé�I�Ή�йԁ�����/�/��O����U�b;n�3�G�����TȮ��I'2Tf�U�WT�3����~X9� =��͔�Ya۳�I�G��s����*��͜B�"��p�>P:t!���&��6rIأ�#�Uo4Aa��cl����Ɲc��S���@�����C�W�]���w}��ɞBgH=h6oS.S.���4A�#Յ[�dbH���M�����ܙ�N�A;�HU�w� �CV�j�������B([���Ǒ�!vd��~H��9x��X鞈\ġJ�J�x���`b����	'��j'5���)v���&���JŸ���]�����k��N�Du}c�Ԅ��du���jMC�_���^�QM#�b�Ɋ��dOܛY ��n*qp��\Ŀǀ[=K ڨ	�����C2�2�S}�����h�n'l����[���G�di_hN�5����& H�#2=7�'�V���L����b�f�eY���R�_P��"۳Y�l)��>B�� <��ż9�У:!��V�JG}����ZuH�t
�����Hy�8�ԵX{_+����̣�����d"	�2��2�K$3�N�2x��E�HД�_@���e�����6X\�+t�^1P� ���̳��'���M�[Y�� ཕ�YB��S-(�������_�R76�zQ�a�Y/`6� �������Oj�~�n��U�"����E�:��W`w���2�ύ��Y+���8��E��ēo�a&Z(,���N'W�TFcg~n
�������1�N=���j[���Y�pd�@���*�h�8���~��g�E�����_GQ�"�7�N�R	�����Z�������2��P ���j3�K��<��$?ʀ�f�Ylf17�lP� �#�ŀ�̮���|��f���u�'h�`�,���؊�Au����"�|R�6Q�S2��t����}>J�4�$�c��نH	Ѹ��(�
	�ELb�)��C5�*蟙�\k��m������~��~G3���nE��J�W/1]Qa�P�M姻_	��C� �
Dј��ə\�I����3}`�I��Y��)���W:��4W�����@mǠS��l�P;���ք�w�͎�� ��h5�	�m�d�V�{ba���_�c�' ��?��b'hDЇ�A��;����Ҙ�*إ�W4��@�dR�(pkյ��Q�/?��S(�{�������lT-l�O��`�@ 8΂tX|h8�#��ǖ@FL{�)u�l2�Q[�*��>���'h_�^0c��\\��L#�G�*w�c���`��mu�	��:��~�%=������u����]Ğ�b���6���|��g��w��~�J���>� �m ��sB
��IM$�L�@�㣨�����bt�DS��v �%+qIj��`:�I��A�rE)�������^�/A���P0f��S/B�HN�L���B�Q��M��_�J�e�)ܗ��kQ��V�v�ݝ���w]U{�e05g�f�c���p9���4��KP����i�&�>G�W>5r�z�mpv$leKՁ���x:'���Џ����m�ⴸ��!��7:E�©�Wa&�5J�o��8���4�D�p��'��&��	hL�ɽ����DF�xҍ�_�R]o$��	��Ɍ����U���@��=�x��?�
ݧ�����}�}��cMTd}`z~p�����5��1~q��hYK�4��.'�6�2CϽ���Ls^\��V�����	�eյ8��U��Md��n�rs��o�w,6��L\m�����.�[��CU?y�|�J�J2�O��m~�ӍBv�@�)���a����@' �nMc˩���Lh��c��� �k�4�Ε��{,q!CCۙ蚑js���c9�/�ᎰX���E��?zԷ�!X��S
�Ĺ�E��h�!��&�P �u�N3�kxz����o�:��;Lx:��Fo�P����rI&d%�ִ��%=��3`Z�@`2\��%PR���f����#����I�H��Zv^|�`�'�^W #�	�;�h��,�յ,`�kN���Y��5��^eC^Ы���*/��_����o�I�X�3�Ӽ"0b�=� �іO�S�dvC+{�y,쓲dU�'���e[`l.���M��P�cQI�q����- ��k
���8�0�+�����=zcD&9i�.mL�)�'�9��^��$�ts��ǫ,[Ȉ�/���p+����`�x�r�ͩa���� .
�~�Nj��~S0�OXw�1���|�V�Z�^��<Y��@�N���56��r�����v�a>�r���T�@yƭi^v�O���԰Q���%��s��'w;B(%��S���r$ǰ��Qm�Ƶ�C*/�#�<Pi���
��|bn��ru��>if��4��J@��!���=
]�F�eP"�����[���p�gU��dgU�݇x�4�Q:�&iP�CM3 ���ݘ��n�`��;B���NѾ�Vy��ǎ�2û�����h&yV�?���=7���.{1,��*GU���Z��z�
��{D7ڂ����s勂���8�Ŭ��j�؀.�p���oH:����9�����~�b�^,�O�ik�̱ʄ^J>�/��o��~;�j�+@�c"S��}6j���bj#텞*<�is��8M�.On���� %E�$2�aJ��*�C��N$�ڙ�h��+
kr�-�����<�M�*;4��2���
��S�qI�W�����۹�>H��
�"��r����*��-e��<�4$U0��I�2A��b������)����Jm����,�m��Ge����v��-�
�M��Ed���W��k�(R}��#;�ț���Q ��o��~a�	��3r)��9�����"M?�6x�pDdi�T×�k�cz��7�H��m<҅�b�L'��9����֚���$����1kO+Y��	��ƄQ0
�@G�F��;	���X�h#��yu�`qu{���w$�*Zظcy�������_I����Q)��]�'l���Ǝޥ���H*�VbN���bC�n^��$f��a��Ohs,�`s���(�X�S�t*d�u��4�7���0���j���[T�x�yqD�f�����_q����l��.��uL6�S���e��GH�,��V7z�W��i�9�0��{�Fzt�w��M�S��b]	'�>4��Ab�Y� 
��W+���E���/���J֤�䤦:g'�2Ќ��<�ePkj}�x�Y��Փ��S�Yc�����a?&��.�	0h¦ryt�mګ�(�f�j-��a��jJ��P%�C ���1l�JS
�S$��47{!n��?�l-';ŹR`\��z)��I���I���yG?���.l�k��h��vIԕ��CU��ل��*�V&3�-�+��5��yI�牠ۑv,V5��a�,��8�C-&n���  �5�ܡ����Q�����1؁��b�s[���Nک��՟���ٌWl�(�]-��[8U�ThЬ�؎�&�?��'}$�L���ma�����MN+H�S��AO,����'�a�_ǫ��o׬!����XE_Hu6�2���V��d���]h��؇���0������,ֿo�BӾ�]l�k񟉠�:o�%�sO�H�\���{j��a�W��=ݲ��x�뛲�sO�Ya:?=
����cu�J� 1T]y���~iV*	H'n�3IK9oF���#1{�P��p�J�3X�e������#>�g��(Z�����CE|�W���b��tU�;D����^J]nq?���������B�W��tm��ą�a��j6�i��7-�m��[�|=�7F@�>�(x�ښޥ����1��M�<� ��u�'[�v�8�ϛE���n�Ԫ�ET��9�d���а���5���z'���LRŞ�!���#l#_���v�h;�<��fK�����\� [u���p�\������Kw��sx�i\���l^ۃ�N��Ӕ�n!�'c����.�������?&���qd*�����9u�*z�QV���_*�4�C�\�eZ�0�K�w�fq'��z#�c*��0���c�'@�j�CS�:8�aQ�돶g���6vjf	�1�F��4C	n�l`���	��ߓ�)@)�ut<��5��7��{�RK����:�:X���.�*O3�jo�s�D�i��ǅ�1��'�+t�~`��u{�����J�zg#��!��i�_
7���7AҠV��3�)�R/�Ot��{����S�^�[��ӧ)���~�N(i�m$�eny$�n]₎�m�;� �,Kvl0cF�/��O�� Տ����ˊ�����Fn����L��)�|��bͣ�z��=�?~[��(�����V,h놠. ��%�kO)J��UU����'k�J�W'�#�6)�y
HX�����؀������QwgA��E!��v3{<�:�7��/�m���k��PU��D�q�7�N�"�g�P��2��lW0�rk�QI�粈lI�yt��I.V��_�%��aM��.��t����m���Ћ�D>k(�[����4uF�bg��j�j2h�R+	42z�e<�_z�8�u���\��VGUh�̬{m͞1��bd�I��as?s|&-���QgхO�o=��6�<���6��r�Sr�_���2-�N��G���
K%:T�R����|����e��{Ř�=z�/���v����61F��^��M�3{Vk��J����ķ�����9�����4�LM�Oޗ@�zy�q���2�C���SO������SE #�������7�ĬC������npS2��耐㶭N���4����w�&"_�k�p�Xץof��I���E0�r� �X�c<~������:�Ur�)bYa�YA)s�ab�km ��BE��iX��#8�۫��|�U�2ޢG��i�欜�I�I)���v�rF�i����4����yg֧,�^iu��"�æ�Kn�*( ���SK�r�����k���C�:LΪ�3'{
����2ClJ��4�O��p�_OP�O~pW܆�G�w��l$�Nw?3l>x*{��4���I�����~a�x�ۘO6wj@:��mEy�$�{�	����27���ϯ�A�jt0U�	�K�:�^�΅mI-�,�Ҙ�m��e�2Q�SI:�oA7�ZU��w���g�.�%J��g ��Ѫ(,rF"��W��s����̽��%A yo����x�p��2�5�MNI4H	qH�����}�$BNo�d6#�*�Mc]u��Q�B9��+gy@/2�"t�Uш��co��;b	��>�%l��3��|c��	 y}�#�Ad�+��#7��YJ��nb*2��0t��Z@�Č��Ź��j�����^�z`�ֽ��,գs����P���N�����v�q�:iz�O!|��e�?ql�LL�r�+\O�<T�t1f��볩u@O�ъ�7���H��o8g�r�����+�f{�i6��ۗyB:"��ȡ�/��N�}�M9�Fz�{@��3����`��$����@��������S+S�'����^�W,����>�q�7Q+�!�@�+��ł���h�yb��{��z����8��g$ax�v��ع�5Η(�|��R���Hh�E�=��yΌp]�J��eJmuY���{%�����s�;�&w��o*�9�P\������!��a��Q
~���b��`N��
��r��@2�+2B��j�C��V�%�X0�#��M�L4�w	�@Sw�cu;��ذ!�8��3C�^��(�\0�whĉ��[�Y�x޽���ߤL�Jk��ė_�T�Opc|uN��3�pvmC�'�ޅ�i�$�'5C2H�Z�b_Hj���F��+Gd�F��V�o|u.�"��c5�r�����k��%��A&_?�s���e|*�`2PnQ:M<]�c�,�0.'0���n1�m�DC�3z�B���I��l��[V;ѭ���-�˛60��jX������W[q��q����QJx��z7�)�.s��s��B���)U�(��a�`J����r���o[�V=b�� �Z������}�K���Df=h�E~���j�L��twhNP��7wr���|��:��rD���PO�x���H��챈JOIG�N8�B���|�I{�F�)��s;�}
�㪝��D/y��U�_]e���}q�L�;I�{~�~0ʚ��HׯG��,���@ED`�����+U�*	۸�L	�Z0.J�z���2a�1 ��Lr�/���WMq��>�vn&�����N��ز7�@_m:*�=A[(�zf@-��c<�zRX�������I @�A�WI�j�%���[�}�FRL�:��[�� e]p�-�*U�Y���9�|T�2���d��x3������=��ig\���E@
�ܖp}��^=��@�����O���2�{�9
��`�P孤�.�>X|h<���)��T�d�ͣ2P�+`2XN�쇞�>�<J3�"�2�U~r�AS���LGCTę�غ��?3���yݰN
��W���~�:fؼ�zxR�+��p|���Z�M��x�DW�a`�% 'l��HJ�%+���`;�Bq�[����!8͡�Ǐ1BNXR�i�Aa�AFk�yf��џ�X�sv @�"�6��0q��(�O2�R�����ff�*_�ց�'���E!tG訹�^u���2�Fi+�2}��ui�!N�{�����iy�(�S�.d��+���R�>�U���^�|[@�%���Y�E������C9)��H8�؀#��	8 	k1� ��
�ӡ6Nδ����T�?�K�o��y�UB���>�xS/\7����*��Á�e�W�2T֒����z�~�>��E
k��~rNMD�)ۛ� � N���鹷����Rx�xK�l�}�7��4��+#�<��-Lu���ꯟ�:E�C��9v�	mM��9����K�\�qh���]��D�NWΣ��
��aM4?%d��Bl���@T���CSt9f�$�aI���՜O�S5��b5����;nu"v��M�-a�������7Bl�����Q���V��j@����4�`R�����+�<�g���.k$�=�`�Q�ɢW�J���T��_͂���) u_0��%.�i��9gIR�K!�%�ӏ)�3��D&Ιh��s3vc{"�,�`"���3�d�����G�:*=����mgע�3ύ��i��Pj�le��5���,��-� F`���0��� �<�%�����h�  �4^{�b���0J��3c'��__�f����*��~c^*7����F_�����9�v֒Jj��]'�Yd�$�H���I����l7]r|�W��J�� �A��8j'�o���jچ��'H�~ �'mϭ�j�����-�����7\2��꺯���a��Hx0/�7"�6�Uо5�+/�e܍<Nމmł���1�S'�A���{�	��hck>�딻�c�qEt>)�ZR�b�Q(����P���_@��h균H� V���q9�b��^3�[�'r�ǃ���Ѡa۴-�-�b�����k��rR�77��H�\�[b��o�=ċn��x���l�������W&u:�;�m)�?èr�ATҥ�\T�=��D�0'_��p[��97WN��Q=	qM,��I�ѵ�ďc�$��q��	>i��o��u��,C��N!�J��Q��0������Y���ѿ����+|3.g�CY)�]A�{�+f��~5e�,�,b0:����5����j�Om���T�v�D�c�L���E�Z�Ə_���W�"���ғ�flR�`X<h?��ފlNI�|X�����~rq�N8t�I9u�o$q�G�@�f�R~JU֒�t���̊�=11�I�-��+���vXK8��;0'�,�'O�oX8C�d��Y�֮�٤:���6�Q�R�0�."$�Q(Ж��)ħ!�|>��B���g�5���j���
 rcF-@��i9 aO�ȳ�Z!ymhd�_ʏ�Tn(����*���Qb�4F�jB�AgSq�j�o"�C��7n\b�v8oJXq_�թJ�(Fu3�u�*=+��7�/dN�fD~�ٴ>����8n,/Y5sI�5("�%�`�h���ŝ��>����{>;-k����/��*;Ne@D�(�9���6��Ϫ��[���4�U�ǣ4�ۻy��V]N	.F�sh�^Fl N<Pt�D­�m�Q��3�M/��Y�GO�̡�̃mB�L8�=׳���W�������F?jcw&D�����#N �=���ܹ���=��[F�~h� �A	�X]o8�M�t�4�.��.��-��煌 !uV(tl���9�{Ql?;�$FJiQ֓wl=�+��n)�D����4�ģ�/���c���\���}$�:5��0D���,��*��~Ԡ���cl��),�.�I<G9O���+7L�zd��!��,��9pt�h'ѷY��;6w�z|��ͷ���2����
�0�U�XVkV�}��o~�������؇q��U��%-��\ !�]<�!����� ��?����.����M��F���A�۱�@���M���U�� �iX���[�O$0�%��h����f���۽�גG�F��.�1�n{?r��Xæ�sIHW؛���Q�����M�אm���%�d��{������Z*9@=���A&��~����������*�?�ɂ5���U�=`��y�R>��O���uw�=ӛ��p)�(+X�Y��n ���� W�a�]�;���,�����H:���G�Qh3Hx�ƙvL������B*�9���^i�����19^�E]�DF\���7ŧ��4�y�
�;6�/��
n��a���9�@Vd:_0~ݫ~�~`�*�f���{0'��K�V�t�5��9t[\�TVT�%��$T����;~ݹ�f8Oe@le-H��hq����+�Z�9��6w)}0��0��L��x^��\465�~��m��W ���%P��ev�=7$r�pHY������UĢz�g��Q����g��F���bY��1��8����Ѯx�����-�S<��}�E�l�����X�n��J�t�q�����TD�@m��R/I0���Ȱ[���}��!K�ܓ�U#yg>GW2V_��M*P|��q&3�J��$�e<\����f �Ȃ�p0@�3I��c�ZE1"��g(K�強Q� ���`�MD�N;�=zVX]�6�f6�Rn2�)���L�߽-˒��*.�,�Z���c��>���D�:��4�NGO�ZǏ�� h�08��ޤ���i��	a�]nƵ����V��,��V/�����������H�CV�b�X��ĕ�0rk:�ð��S��s�+�H:ol �ۊ����c��V����4W�K*5���ā%h��̲f��cG8�-�)��ПB���pk4�@���(��+�T�~ �Ղr���`�T�!�0����l6���щ�''d��8�L���F��Ί��O��mH�/�r�of��q�q�����`Tەff��zCǬ��x�8-��'/�����M1���L�;-U'�|��@��2�g��a����G�*��:qh$�LH�F�1��M&�Œ����%�8��a4B��=���:��\�2 �@W}Vh H| ��k�I�<�� ��z���oU�e��0c�q4�]c�Z��ޘԷ8B ����\����Å�屼����/���ܣ��b��l��6DN �<�$�5X�}��)U:+�dH�Qo����Ʒ��r�@�1�@փu}�5A�'(��|.ᗺUfF���AVdf���ag钔6��4��K��v�Zxs�{�/�fC	+#�uQm�1�O�(��I�R�u��x�,L�|>��ܝzN�m9ϫ�#�H�K /&2l.�2*�q+�D�~���
k.�\�X'��e0��ԃ-�~=�:��?��M7�G�SN�e7��3��n=f�.���9������kA>��\�`�dڄ��SV�C��~Ǎ�Ϥ!ƈlAf���^�P�М�CW�%�uܮ��?����g���uC�D�V�S�U�]�٧�F�d����S?��Ƨvɹ���`ޯ��G�%nI�{���k�h�rd],��wq��ر�H�c��\-�|�lj0SŚ;m(�xg���h_�2q��o��I��۫����ϫ�>͎B�]�m����f%��R�خ(�^���EfLP���=�����G�&��bX d���s`#h>���܇拦mR�X̿R��I�$w+Kl�Y�7�9cx��S*�ͣ���r�:%Z��Uâ�4�/K�� zmf?��!27yt�Cʨ����m���S W��?���wW_�k��`�,�� �Y1`Bj�K���Q�� ��ݳ҃L��c���sx���l9� aeyT��OF�9����(>��턡�N���~T�L�z��2%���_�SW�!x0E0��<�]�F���&c�ª[�G��Ҽ����%��	C<�,�����&*_?%7�G=�Vv��Nm�����-��)�"V���qz�mj���#�1;����i߼3�Wǉ=%e��"��sm[e�°
v�@���G.ܙ<B�XܠoA��V枙���8n%+�.���<�jz�nBs�7�����$�̆#�zl���e�MXU��|��Ku'��܎��2
��S���U/??)6����^���@BO�= 2��C1�U��ǯ_�K1㸇�M��ŹM���+t��8� �a%�T�����&���mGnA #:�3C�4~�s�9I�˿oԑ�
�߯�d]��G��z㼇I��<Z!��TAQ_R%��F�?v)��z\a�!⨀7*��sgA)8���(X�>�2�����ɐP>����?8A��9u^s9�xv%�7$��c�}���@�#<"N��z�0���H�[1|_�~<y��8k��i	3Yu+/ikd5+��e/e��O������.��m�Z8�u�|��9�V��Q��eY�ਠ�9�{�+����|�SW��{�m�@R���_I<0�}�l-�@<�UR�������bdqQ(5�;nn��V�!��:���+��9�,>�Z�Q���)�MEX��xL�IY�o�H����qT7b_*�V��:�Pyoȟ3q�1C�!���`������/=5�1C�36�m�3�H;��r�G��9�+��XZP��/a��7'�a"�I2��h��ӥ!;�e�����"]�+K�Te3ܠ��J��|)	|�0�12���0*gƅL�E��|h�[*{�Cv�����ϒ\���-]�h���R�8�&���K�S�Rt�B�4];��Q`bN���*�������úf��:G�rh�D�R%�Hb�������ț�e�������χ��p;�*�s��Ue���/%ũ��8���6Ԕ�r���'Lt�ήt��W��\�l��b�#d�6I�L�F�a�E����֥X���|�^�WG5�D�Q%W�x�P��$�Lq�K�mz�|�dW'���g�P�7#��)�v���Nĥu�.4wեM��l����TL]�
���&�.��Ep�c��_.p������1�7�܅2�cY��攰"��C�� 3ю� 6_J�M���U�C���|wM&��y(O-�U��)�Qp��TJ'&�6z�J�����3�`d��7S��	ĕ��ӫ��b��9m�P��F0�J�g8x��βO��"���OAF�����:bz�ഄF �������⹮R��^`Ͷ)c���i��d<q��$�`\�-��Z��]���<3.ޘ������0���8*OV{+/�*�: ��\��{3b�u���{�uz����m�?l*��HΠ@�K���+/��{jj�J�cF��-aBR�/�������2/!�x�@p#�-�"s�{���F�QE�)�RZۺ��:���8x�h��Bs��+lM����I��˨�-�W���`'E������7����)0�������^�H�xe�b���G옋���~(&_#�u����K�2uC�i�2\ԋ����t
a9X+�p`Q�4Q�w��  �i�D5KzJCn3Q���wev�hގ�d��C�ݠL�}��M2����?�&<C�Jq��%KO�,9�yey{Ba���M�$/It'b�/���D�&to���:�Aa��E�r�T�1@��d�j���7)Ǿ�]Y�r&m6�(w �,�}��=�u5U��ɾ(�i�Je��v�h�\��IFq�6�&���*0��xk�_��֎����%�`J�o��&��CsZ�
k�Ŷ}�3����<8��/���)�d�X�Ǣv|j��aa����ْs/,�C�;�1%�MA��.�v����lf�l=+���VOc�)���U���t���<�;��[�����/]�ʶ�/0��]d�:%U�Tu"�Q���vu�6��5�4Ľ�����������uLpz�>+�)���D
���|` �A�]t�(w\{.E�p�/��V�9�����6N�J®�#�'Tߧ��h�׶x��+6��m0Zk�u�t��nҾ��8H�*���5�F�t*���Q }j�d� ��%n�ߓ[;��<�d!Տ�3,��1��!��~=)�ZvԽ-M��VQ�]�*�N��8Hi�l�-��-���-T`
���٣�`���b���ෑ��0�޸����e��>�p6֤1(K����h�����Ҷ�I�Wq��0�Ӆy�n��1+f��[\�/s&����N���)�c`�E����P���N�qK�7��T�$�g�]��(���R�u���עq����'�l��US��JJꬠ�V��9(b�R ���r ��`ؾHh3#�$�+�F�X�׺�"�J2Ĕd��#������si��˳��3]P'gP��}�.��m`��i�TT7R�r�dBps�V��d/Pm��#�_YW��h�"�U^�)��|�8PB��>P����޺�z�����
��+6�nBr%����^�W��̷n�6�c�n2N�ٌ�θ���r�x��<]��À"�K��CM���_��������Y�I����k�ќ�ٞȍ_,�zx�<n��Ibb�ѳ�1`�k�SS���'�'�kk�U�*�%��k��´At��\~D������� ��m�j�9M�ܸ��V*d�-ѻ�͆h�g���~����B��Y�}s��H�����c��i2=U���Qy�W(	a	�'���}?�i��|�����rX5t�\lK��mD�7��;F�F�5Yl�a'`�깫�ݱ�������#c���M��[��3"���
O��'%Y��X^}T<���	����rgz�fs|	�eΎ����fAɸ����A���ӑ0��S�, ���:�_y��_����%�|{۳$C�	����!�������A�W�f[�dmRB��NN�9nU��K�u�Z^T o7��Ǖ��1�S厼�/
�/V
�1��6x� ���A��s �!f�xwY_D��:K�Ͳ��`�n�Hi�3���> oG�~�oخ�G���N�r�A�xj��5f�t�2a���6a�*`Y&hF�ʤ��\���Q�Nm$£"A�D_g�A��i�\~r�F?N#`�k9ȏpס�Rb	�&�MUXh��!�W��k^�Li�+{���pT8&(�n��v�� v��H��듥|J�m��U؍��xq�J�K���j��?O6��;D�h�O`��)z���[.��e A5bc�GG;Oyϳ�i����=���P_'3�����U�-X����3��p,���~���&����TL�2��^ȺY��&�������i�D��>�����Z1պJW�& �ň�x�^M9���5$jݚ�\�X��3o$���-b���\F���"�w��c�J:�<�%�I1+�-~��3p�.����Vf�$�:P/&�DEr�P�+����{H��ʎJ�෵x_���^~,N?�Vu1��?��"  V��ԝ,Zxf���%��2m�Y��f�r��WN�,���E�uܾXU�.iAL����J�埽i{�LU�5����#���*����z��9��u�ROs�hEv��S�V��:����%��/Ky���!&�)����z��sI�=%��
|4�ElBqM3�p�L_7�K>�uɕgk�sZ�2f�Y��`��1�_+�ӌ�o=[����z�~3ɯ�b&���Yt�fM�I���[�g����ߥt�'�f�w��7�F0���/_��o5�����كW�z3��j��i歙�5�p�m؝���v�e�T�� $�4��~�J�{��}��q�<�E��ݺ��K�~�[
��i5��JJ�����%� ���5�[}/)q�*�] J��W�&3�e����Ξ����Y���^1C`�(b��=�o�>����+�*e�⠰��������=��nQN�YE]tF �ݼr�������/�T��G�A���֋���kFo�"&ub�f��2H���A\�>�끻jp5���'	�ߺ�~��?;ԏ(����Ɂ��[U#�꣩+c�^y��A�69��18��F���$&��WhO����q�M	�lԾ~�����Q��Q���7٢�i��_^bӪ*����������_���Q\/C�E�kV՜���4�`R�%o�����)��0n�.rW�*It��W�F�xh�n�>�G�<�����������O��q'+�cE�+��"4t��[�B��Y�P�YU���Џ���SA��5��'D��}˩�n��&��Qڔdw��u~�*#����*A���㒽h"�os�`�@�S�����|X���o���c�+e�Y'�b�o�*��ʡu!6���H�������.7_�zy嶇�+�#䢊ց�L�(�d �b%��Ŝ��(�}�kH�����,z*t}P�jM����~1�*>=�{��bE���ú�|n���d��T�!�oO7��'�k��k ��}1�W2�?�)��3�,�;�����>O)C��M���-��m��<^ol�uqvx���]�i���K�q�X�XZ�ܗ��S��0vjoo1\b�M~+D�W�z9�"���H����0]İ�:o1%�Q @��I��]�MK~n���s1�[�4�?��_]ګ^��'
������`޳�1�˶�6B��\.ݺ�$��J!؀֩��qG.����m�aI=" �о÷G! |(3h�ۊmة�_�K-2w���:	Q�}�$�6,Q�\K�mO�G������P�6WtY2�'y	�P�����A���s5��T�*��J;��a���gƅ.>�mu5�a��%��F��6y[HK�&Y0�Q�W�j5cȍ����c9g%)��k����1�0��c[�sףy.�#{C���V�R�$����"��y���K��֑���
�n�[��������B"��.��"U�;�Z}�BM�/@�Χ�w��g�σ�s�^.~5au�`Ql9���b<B:;�'G�7�]�KQ�Z+H2_�o�ܣ�=C寏o*�&�b -no�I�ow��j�l��s7���ߢ�}�BD|m`�_����א�����EDP��LNG�IcJ�1摺��+sp�SשD=�J������~�4}�{rɘ0�1��mhP���'˪�L9���n$���fD_n �����'�ny�I��(@�+�7�ަ?����o#6�������{0�L��n&!���/>�N�;%�=�����kP��}%�I�h�3t�����0�V��^�E�L�kg���[UM4���=��Z�;����
��iU�"}Oʸ�I�d��6�r�'��+�nꂩ8�z���Յ�ᙫ�|�|�Т>��Fx����)�?<�$�P���~&�}9}w�Q�b!��TP�㔃s)���Rhg�kS��`���b�ɱX:�F�pY��@j�4�Ճ�P&���66���3_���˟Lբ"%��$�Rr�\��	5�g���J�A�E�]���ZU���W�Jj߿m�Sx��[�6�R
�#۬�B� �\%z�{�rK6_ʕk�!�/���%�I˛��~�!�<���_���a�Qy��gR��:���os] ��)�LMy��5�:) za	Gd_Go4�VU��G:dG�D�^WnV�H?ڡ�C�u���Gl�ͨ��V+V�^�V`����2�w�W3���z��|��X�!����S������׳hn��L������x����l�J����GN�����Ļ�c�r����3gQ'wk^( ��<°g�/��*6��.y^58��'y����g� q	?�@z"��l����b��2d(�gBp��d`
S���ooc������gM&�s2ճ=��iwZŉf�	���/Ǆ�K3kI}!�@�����tF"�U���~2�n<.���M2���R ʁ��!��ǲ�c���I��������L�j3���.׸��3n����oGw�v�Q����qQ�}� )���-"��Ѩ
iz��%���8�Ξ���N3��n$�5�F���U����n��R�+8�8"��u�71`4����i#zT�S��F�AZ߽
�-^�Qiy�"�W�'�Q��vq>��i�'٫�Î�����]�d@d*,�î;�X�����ɽ�Bjf�G/B��Y�/4U͙��Q��(J��A�a���'�8�/�c�WM���]��\�KX��G� h�7)�
Mw �C19��<_b;��MP�p` �ak�A�!�8~sK���#W��/fI����:"��XI�!�aA�6�����lމba}TKIcr����{��Ϗpm�\̨z�J�(��VJ�<Qk1~�Ay[{��B�]��q�v"O_;�����G=W��!Ih��(c&ہ��ڰ}(��+h5v�5%,�ل�M!��kJ[&�\i<�������d�~#�z��?S��b���n&���<��y��_��8E}	�V���i�/Bg���P'1�/ػj��M#�F�>�G�/xJB�4�b���V1�? =�Z\�ɼ��K�|4��ʈ�c@�7����3��w���X �mRL�	|i���u��h�X�n<	�u&�5�RV{�����SAa,�5�L����==r�鑄mrg��g%��ݑx�,U:��7�"^�İ���W�[
���)����P�%�����j�2�������yGi�`�WjC�b��FK7�[��]�f?�_��<�?�ݝ����4E�<�S����1������$��Uj�V f݊eR��7Ɇ���r�Y46�}�2�f|���T�Ł��G�^_�*?icQss�LŒ��~�^��H���gxK�(I��3�1��}�3�%�w#×�����o0���D	MpѬ�[��t ����-�(eMV��Ps��7N|@w�/Ȥ�Q����70�XvK���w�-e�|��>�$��,l������.���z�*7��g�"R��:���F�'}[��X�-e��$Y�t��cظQGz�֦nh��[�C�y�>���K�%Fq)6�j��&�a7�8�y���A���z���e����H_|�r#�6�RG�&�_���H��������"��q�t���>U�|�S_ ��T'8�'Y��x5v�D��A�R�J�7W��K�0���q_5.9�@�0=������SIcrr.�,o�SY�}&?��6Y[3c�Z����"(�w�*,�~�&L�)+�{��7�`�lE��9��n����W 1y~��f[XٽV��FQO��<�9�����>�����&��{�$0(פֿX7�.cf[/;��r��|̨�=��������s��V#��� -�D�*��񛈽���8���-M�06�����H*0���h\�`���/�K��~dђ��B�Z���+F�k��1���Y���7R�pن�������] Zo-h�kCØ4��Z���00�XU�T/��ݸJ+IR>A���#��������=(��-���/�W�U�jekO�������NN�6�Z4��q��^db��A����8��� 0bB���O��Z��a�Hm��G���`�<o^����[&6�R�]|���>�spT�L�]w~"X��T���ݽ��a�Oe�0ɦd6@�i�<O���L�T`{/�V�<R|c���iP�Ċ�Wo՟{ �\�JՅ�!� U �c.���K	��I��ܵ*��!�X���*̷v�</�DΤ/�sw�>�ʵԆ�x�
HJ����M釸�:*�^���r.��j�oe�?���r�vW��jv�Q��?���Ƀ���h��֕i�P5�[�4A����Ⱦ1��qq�D���U<XmN�H���Al���3�.[� �_drD����xoF�6uW(�s��LM\'+���V��	B!ZVs�Ʃ���>r�u�Y��m��N6�n�Mh6�64�!:D'��^�����T1˫ՄJ�N����+��t��.������' ��,�1pϯ��ƮJ @=}2�,����C5D����!�~��^<�2�=�+��SD٦Ģ�)�=������lЯF6��	��ia*�2È�f^>y�+�L�-�C���O*ծ_IT�]<���4�����u�M��]��:���U2�i��9D�݅F��́B�Hٙ�z���Yc���a��lb6�!/h���3^r�S�0k^���b��N򪏯|�xc{輓��Q�A����V*�1�!p��nx�PD%ӜQ}ѫl.`ܡ;��iM5������� �ƺ&A�i���)/�	�)�j�>�:�X��I��*���8��PlP>;�k�����g6[�I�/:�4��F~�O�U�@�kZ��t*gd�Ռ��(����6�b �	���E����g���M�r�8-�6�+_�e�s�r�R,�t�I�=���s��]��,*0Ū��7�?̦'�Q�>k�a�;ؾ�O��%1X5���q��b��pk�D|q{
w;�Dg�1��#��||���X墤�ɋ�e��?�T¤_�7/�f���L6�^�V�<L˽	�qb[y�����gs���R�e�;��	�Ȕ�4YN�.��T��75�Z�Z]�U�QcSC�-st�Z�(�|����s:�����A��jX瑬>r�����4�HO��nɽ��D�Þf_j{0%���|� .v�#l���ΞP_�s�A�I܊}4���m��ش�l���Э;����i��UE�BC���;l'+A�.���	ȸ�k�%\b�D��ȭ��k���O^@��+ys���p�����(2��c��Bj"�Yóf��M��.=�;N�5����oΥ,ze�<Ÿe�v��7��SB��|�,�Fv4�҆�+s���@u�v��ǹ+?�?��>+��c*��n�f��28ٟ�P��70B�Q�9�Z�p55����s3R�r�&�զ0"�*Q�Z�d>0�P��1l����|U���w�p��w�3�=o��?����b?��B �bmCJ��Q�YRm�ւ"C�2��S�@��_Tz o��p��lr�O�Ǚ-
m%��W	���	�AJ���J���0�@�� O�~��ʭn}��\!R vʤMy��gKIL��ux�$	���$��)&ー.�� �0�"u���F+��[���F�7Gx�\��0�&�*�	�t���"˃3o�����*:��AE��E���NEfob��E_�OV$*������D����P���nr6��m}�#���I��U ��V����i������,8��Y�\~�.��-зxU��b<t�ƻ���[����8�W�pU���M\���bʙ�6�	���s�W�Έ��LĹ��$~|��f�y��p�̹I���У�dt 3!JJ,>b��T՞�:�+�'^�z����tq��� B0����:�<g--|��C('I�PaƩ�&�%�V��f�Yr�xE11�43��=G�BIj��F���٭�yWq+�2�y/B���j�ﻆl�
#0����j�O�.��J�ү^�]+�䌿���$�b<�+�]�����P���8�V�����X��Ǫ�JnIʹ��;ן]aS�� ��q���[�+��`.�n���k�c�-�{u"$8�t�'g�|!s0�%����7��N�m�������
�1����WЈlQ��s�@�34߫�Bg	�W~3����X��FPˊ`]E
`�Ax���֖�X������]���6�6MZ�⌇&�U�ʑ��ɋ
�H�ʑ]l���P!iq��i�o�ⳮ�(����Ft�>d��#�F,}��cqw�u�ؓS�z�҇ B��޹;����U,�&�s��̤򯼕Y�E������v�g�cJ��?�>�g�E�H�rUƷe��"�JkI��>VP~���?ۛ?�[HG�-���bx�u����	{�pg��X�K���?ŌE�����n�ă}�)N_��x�H�����լk��1�c)�y~Z��G�C��Z� ^�!q1o����!�=J7�'�P-7�a���ݳ
np�5c�����!tʆ�O���%�$0��Ck�[�o�4޷���fϘML�)F(0����My��ym�x'�M����gTs|��%KvZm�`�1eL֌T�<~
�!e��U ��S�gǰ���Eyp�7=!|�0�o��*���<��_��g�1�U[��~���T�JG��֪�)m9�W�2j�b��x=�*n�?�n�Tj���aF��#���FX (��o�u�f<����5dڥH�%� �}x��H��F����9�Y�� �ǂ���u�F˷�����ݱ)���t~^����b����*[/IUc��5�d܊�9�
)b����DMA-W��YkcQ��(�.n9�U8y:�Pr��d$(�����#8�|78��PA����h��gi��/�R&�M}���!S���C�>bD�5�M��5|z	b\��V�>�U���UU^��0���U��n�Bg��u��t$�����j��Z�.�P���C/V��Mn�⾡8�{�����1�³����jf`'�^@�ъ�o�^������)kD����cYJY�]�շ*��.��$��fn�7��tCm=��M�_����+>8כ�����]�ƌa�h<>G�5�'�7J��Yl�m�t�Gy�C��VT�6���
�w��F�B�H{�v���������R�.�ғ�r����}Mv�z�l*�qt�;���Tk�$w��F��ú�]���0���S�ʄ���o^VJ�OC,����<�SAXd�����J ><�m4�L��KE!
Yyl.vCM�q�2{�o�.j�f˒�%�Ʀ�Rɓ>#�_��,�Yd=�p
k��c��zQ�y���(U��������c&_)zn�[�p-x��+�۠+����ϋǁ�6�#���Џ�] c܎�}��\���s6�v�
�n�4�'?��F-�b�d��<< �x���B�t9x�����*�"*��tUV�
�	$�龯�����2p�5R�Pu�<��7��!�fȄ�ؠy�[}Z��B�$O����?1�깰����� .�P1i��23�B��:�.��`X?���.��˛X7��E���g��BoOCp�e�oӕ�Jy̛Q���m�~1̼���`���1t���|��So��j8�4��uԒ�q����?��\��Ɍ3f��np/�[2r��Л
��M�7:/�$��Ƽ �G�������2�g�jf=��(-W.�O�36� ~�8���6�$(A��M��sU�
/�Q�̲NL��o�P��"�vp����
��RP�������$���k�;����n�׼����`�}�r z_S�W�x�����%���Liz�`�f��Y�y}��5�b� 
�ڽ�D �%��CGm�9�>>�?�m_�Yl���8On'���.�d��LN�QK���UurT$}���0�~�Q���H�3e��vH�7�Mtv�(0��]�n�p�GUx�	x_�T,��.�5=�ʪTw�6�4m��mn	����i�0J1�4��lj>���Lz�Ki��RK�P%s�(�f)^;4��Uu�ᜲ��v�;re��2�)�??�����l	�LxS�����ʓ!�Zqܷ�4`Տ(x������@E��׼��Dx���)�G?{�8EZ�J�9YtX�Zb�Tc�K2ӞÞ^�]�Q�LvU�ʹ?fӇ�؇�O�,2-�~a�%ǖd/TAN,G!��ĭS�lj93����$X��X5��$p܊-FS4Y^惆�hM�(5JdMr�,S^�){o��t�*��S���+x��9����p��t(�n���?��F1��	�(��z<df�;�aR��6:Ϭq�v�8�D�9)��G]�>O�{��Z هT��;���(��h�=�V�hLt6_�����=�A�>�g�p�oEl4�*ϻ,o��~cI���DV|�?;���yY���L�&��ms�(���Ō+Y��=�vi�<?`RMLل���kC���yO��מ��yE�j��8�N]�J1�\!ʟc��VkWJ�"�f�f(��I��\d�p�G��V�A����]A@�|�{��YjS��p�c�e��l!)���L?Հ�B�m�|pRSʊe����T&N�=�v/��H��W�D�^E�w�s)`?��6��̭x��Y�NF��(��~�:u;��|����-�E�s��Zޭdy��N;��O/���ګ�>��}!�/�q%R�f��E��R�ǓUҼ��OH��<��f���?��_�ko�Gʝi'��S}e��#s����q�=��C����T��u��AReC����_Я��91�
̂x�&Pw�]�2[
�[X� 	.�v�Np���B����T��t��B����z|�b��\�c�p�L�� �+�jw8BWES��}�YtgNf;1C�bXӾ�����!����IMT��h�"&�ra������
8Ģ4��bR���{��@� �q�]��6�������z�L��� jզ�?C\�e�4�j��Љ��cS���$m�hV�l�B��JR|+;6P�L��~�;͉���D��g*q�@�:�f��>>8�N�V俋�7�)�Qr2K���U�	(��C E�z���a嗭�ы1+�J�c@���vSu�����r}���$�����3�@F�P��ť�;*��'�s�T0�K�S3��	$�6�"��b1�P������uʺ�]���և?du."8��(����$���j��+����Ci���}3�3��ԓ���0�$A�1{$C��Y�#����*�k�]�tW$*%_��x|ѣ��yX��i��~��<�Ȇ���ysԲ]#M�E��]o�7/A�^L'�Z':E>v���s�)��f��Pc멀��>��Yo���2���[�Õ9v4wp9ׂӣ1;rP�J^D/۾QS�^��+��	�� 5:�P�����c�!�J �t,#�]n+=2K�_e/�Z�w9����"cƎ˵=Tr����|/�6�uC�:�d±��Š��l�����A�����8�M z��[w)��|��d�����)�mlcyL��_F{?u�^:$�!�a���N���j��Y_w�˭�u�ϵ��U-('����6����b�!R8Ҹ�Hر�p��s���8�T�2�;�f^Z�u�������K4����ͯ&�m�o��D	�,��C�d|��]��Q��z�/���q��$T!��|��Q���P����E��2󙁉����"Ǘ!�]-���Sy'B�?�����5f�� +�>�i�y.㜓6�5�n�p��>����T����ӗ�$�[�+�Aߴ�5զ8^.ȕ����.�dj��n\���q��)6<���5�9L�0�����mB��O�Iц@e��P*}O`& w�kkq g�fu�O=0�( ��/_Jd/)w7� �c�z/�lL�L��_����G�y�r���sw;�Ӵ���`���	��3/����T�������r3X�|�{�
r4��I���<�Lײopjrh<��^����7�Q��T�%�1�WE�������m�����(x5�yu+E�/��l�N�k8����i�&
,�N��{'���c���Ns*�QJ��� )~�B��	,�%�J�٘�K�q}�K���|i�1�w����B�rM�=�(����H���G�O������*��EǞ�����R�6�q����E`�Q�L���PS�G=]�w�<8S�k��:%����!�Y�^�B�FQ�{z� �K$�Ň�ך୕�x��|��']
tE��5��E$L��M���1�	k����4�:oo�%���L-,:��w�R�b�3������S3�	���K�v�"ްKϫ]ĭ� NBX���>������ꈠ��5��5i)L3�]6��4m���]�k�T��'u"��WZ�w< b�����@�P��l�x��:BF�w�i����*��@P�A��'<�b>�Φ�q���rw�>�!�9����X4>>K)��ɇ10��,j5r,��:�Ey � r3�qp����>��6&�I��<�ό�=̝K�p���W���Rb#�4y̼�H�W}�uޅ�L�海��5�@�(���� ��N\��cڪ����ūz1����=��V�����?S*x�&$j��@�ʀPA�CU��tx����e��Z�-�(���ѽ�<�G�;hEL��g�I|M�R�0"�i3Lcݧs���a_�,俣6��'�첅N�ƒ��=@WG�Xҧ�k�=<���k� �[��m��du�s�i�U}ԍ<�G(����4�&P�[�~kk�j�q���q��`��;�j1�׮��}�D�5Յ��^�e�G�Oׇs
�������Y=]J�N�(�Y\���.t��(��$�^m'���v~\궫ߵ2������\�r�|o��h�b�*j�ptAI,�J)�2�D��}C4>	�
��M�a�I*���p5�z.�?G��Cn��0�N� �IU�����β0ã��᝱�"<��G���kĜ�ap���jU�;�j�+��>��]	z�x#�������g.3E�<ݍ��R��P�T־�\F���_�����!\�?�X���2�z%�� �ǲ8(n�;�=$���Sѹ��,�k���+h(8��Z��i),�<��P7�_�Mw.~<�^�WP��r�]���D6d�g�����%/w�>�\@zH��fU�N��[Zg�$@�Sw��� �D�V{)p��&ac���9���䖾v���[/�4E��pkw�1�ׂ�u�1���7ӎA�MX�ӊԚ�bb����8��ޅ��ڶ Z��v�pzJler[S\��gP��E�@��֋;���a����B�|��F=8�d�UV��m�Z�<3"�f�獐���:�c��Z�u���e�܄l�
�������o����eDt�
Kb�V��F�(��E_���-1S�Pe�n�P�-��8,�p�xҤ����Z����%H!�ꕸh��
�0>V-(��O_���pU�$��uF'*]N�.�T,ܜ��p�=%6�ٵ��R�%�y�`}����z��U��F�wd��x���m���P���Ɯa~Npp��IL&���S��~��-��׎\���LP�XΑc��X���w��qmyy$tL�W�
�I�EB`8y%uL� _f��c��n'��^�8�b��.?��wH��> ��~ ,w叜-p67G�$n��gCT�]����#�*G?NVT��YAo\�u)�
�hP;��
�ƇC5~/f�� �ra��
r(�1K�븻t�9� ��̺@u��� i��R���O�,z:�W\��ⷦ���Z�}˪�D�v��a���E\�9�1��?� �-}z\'w�ll����l��ѭ�C���礚�r�����݂��I����c\[�/�{?&&6^^��M�Ij��֘B2���r����jzz>�����f���Ճ���F͂��j�����dl0JTY�:i�$�Ū]2��:�eUJ��U��0�l�2m��y���*��3�?�i�j�WZ+�dZN�ɦNܦ�&�@��2��.!Qʒ�XwV2	��R��a%���Tx��+`n��9N�V�y��Żv�]g)��}�(׊����6}��ȇ3 ����7�Y�?f��)8""تr�:߳�4۷��1$� �h��	!X��6���\��	�
!q��M����QV6
�/���~0�w{m��q�6��VJN�T+���q�;��J���YP�v|b2�N�'+�M���7&o��p��'=���L����n�twf��	{��}�b3d6�kk�Kr����1��1�E�k3@��z���K�l�(�s��77��(<,�i�B�Z�o��)k��ş��X�����10Q���������9�x�F!;��*'���Pe�����SS��K�`�ep>�Wqj�I���7�.��X�_'�DC�L����`H�W�b?p�h����Kb�9MYt����"�}vV��w�)y�/�T�\�0�'�}g�A����$3���a����c�TO�*7E����o�7fp��s*\���kv�DטV� h� e���V���0U��T;�+��_�$��W͕�����!�6��Ro��D��ےVxH��{Z��Q�3�qx�����+��d}�eEʹ�Wt�Q������O�Z�e!�i�U�<Oy�[������uƑ�Q.�zUBIMNևp��X;V�d?
��/��r1�23���C���KZ�0���&�*=���`j���1����Sl������J�0�EJɒ��׾Q{�P#�RAb�b��95F�2�}��8��'e4N�q2�8Md����oa]
�gR4�00R���n�yI���mW����1Z��LИ"^
�u�uϼ���c�D��3_� `�=��I���矅;� ���	���^Q&Ln���}^&J�&^p	�#�e(Z�SvJ�]ncݫ���A��_{p���Q�1Kb��-Y�D�&>!xm\>�x��Қgӷ9�@�`�/�Y-�+���~�~.oʄm�H�eĂ]����ߝ�2�c
��T��6w��5�{�|���2T�.(��O٨џ���W}$���o�\�ϔ����y�����c�"D*��pp�= 
ϸ=D��-�I�_��ے>�(b=��F��%�9 `s)�[.u`Y�]+�K$a�0��d��`Zv���K��`�`/��4��̔�L����f��~�g��xc���M�R�0c�WeV,�cO/��D=o��1�)0R�㟨(���Jl�C��tL�q�����p�����B1��a.Y���P?s뺿A��3������R,�,�{ݢj��~7�p�kWd�Z��8���(�½N���;�Vfb�LN}R�!��ۮ��Mt"�N���=�TڡH���T��;�����*
�/��A���������Fݷ�{�%|����fdt>�E��&8=�r@`Km��������蹏"ya1�1)#�N{o�ʦѪ^�Q��,�y���n�qs��K:p\ƽ�c���ܻ�� �B�����:�""&�2�Q���:���e�)�w�C��$y����0 ���p�Z`�KPH����?{��:���A���-�og�Bi}��x4������I�?�����F?j� g�%��� E؜�U�x����(��T����k2��x�<�k����z��I4*�Cq��D[VN!��|������{��|@��p�<�r�����6�?�(���G0,2�J�n�j�A��pkbj�+^�2d� E���k�\�j�d�Ë�^��؛�����8���#FH��2���]�y��,�����DI0�Bd�\�i����J��Pl���2S���PQ�"ضuw�����K���($���L���xEzx���^�
�?z�o1q��<�?m���n�c^��8�G�Ì�L�p�$��v+��=J��+h���)KU�D�u���C�j��9ͦ��D[=妿�fAp��Z�Ӱ��Y�u�h�*]��|�f�(,�������ڻbK�)G�s�\M�r���{����P��Z�<�΃i?� D�q��f�h�����z����*^�jB:.��\8`�K�3���v��'�C�_�.�RqA���t\�'� bP�I
AG�.���<�\���/���k��d����4F�hi�/�/����Y�]�=oA���Z��i�b:nK��t��i�Wz����z��ٴ_�N
!�$��"�Q+M���{��t	�O��}?'��m�8����3t>[�spjTJ��9W��Qp�&m�a	�mG}��,���?UƯY��7H���x�@&�y�D6{}���*����� $WڌR�6�����m_�.��~�U\N�򢰽�{�����H�.��2�D��ݜ�T��8���.ZOD���)2��r�o|���6�י�}ʋ�f���6J�� �����6@���5��,f����Z���I����١�9<!`�7/A�6'��FHQ�c#��Ϫ��~���	uW0��V:;�
6�C���Ŋ78�M�{��#w4K��@NA���uP�����mGG�kyz� 5�퇻��@	R��»���m�#����G4�����-o$���
��w�,�+{3p�p�/�'���H��ʡ���bB��>�:�'HpIjz�(���ۨ�yPur�����Fo0�|r1�h�f{s��s,��G
�x>w���.W�
h9~ύϣ�9��)<6ޡ�	��'�|w5/��.�����
���@f���F�Gt��'�!�E����gξ�O�}�.�����nmI�����E�E���s�T*�U<�N������˖����E�.�BXM�$��7�i(���Y���uJ�a�%W,���
#���u���!�f�b�A_�['l�Bx� ��/�lȾ��hy.��Ɂ�DT�6�k$��S��6�٬?N��Rݫk�^���٪��_�ޠa�A���_ޘ��,�M�=��v��j�X�!�?��_ �Y5ƍ�����H�N��,��d�n� ���X���˦�|	hg$(����of��O�fÁ��!��%/��Gq��鐁d3�M�(~����a������8pS���_��n(.�u�x�/�[(�J
���.(��<��P�@��@b�g��P��λK���Rq0 �DRX,��s6�,�[S�NCL_ =w��ޖg��h��m�Q�-+�rX��ca�D�a�*�'��Y̬<�;$�V ��7�h��Ȧ~�M�"''*/.ۑRy�d�-����2s��#y@XG�8)���P�o��F�;�u�wǎ螺��T�AM&�ܦ"?�v��\g�(��gd͎���֮�!��l��2_ ����!5�+B�����ѨT�1�"�wח��8D%����q�΁�־��
�qNZ-lG�5��?���7���qB�I1�
�½����&�T��KBr��� �/j^힨ʫN���6�H����h��;k�E��Q�������kG72a��S[��	�������	z+L��(s�\��WUPR�>;1R�I���dB���ڷ���S��SC��I�Xy��p엾���]u�8~��)�Ko\��3�̙��Y��� B>�1������!����z��M{·\�ծ�&;���+�+�Uu1K�?�	Tc�B��[��BJ
6!ڴ�{H�<�d�l�)s:EC���EY#]�&�����_�}�,wc-�v�Cy~�������.{a�N���TN�S�!�O��fa�x��ԽF�wc�C��M�Xq6k� ��d�������ɪ&d#���4�i���J,�M��I����j1���x�-4�w�$�H-I��PĿ/����OA5���2�Qaq�c~��68#,)?\�E�v�;.�@�}2�I5��d/AI�vy.�.l�����t2*��J ��<d�D�L �?�ځ���H����k�b�ۢ  k�����l��L'ȁ�&�1�����o ��v:w�\�����*!������������o���W�i���d�F��d��8��p��� ���o��k��b�0yv��懳3b2�NrWz2����#��p�������2]��{�K�綁υ@ �m�n�=���Ld��G^G�T;�&�$���+�9���j͕V�P{�b��ηu�(�K��0�@���t	���|[k�-��?�eZ�)Eլ� bW�0"p�R�3b�Ԑ��`�nו��V%N�M�8=���=�#[b�o/YxF�R��	%C�U(� �A��$g����r�d������ 3���o��E��2'�rZ؟��c��D��'��-�p��ቀ�t%Ơ����'vh�|T�QE����	D��mPS��U��̕^_��R`�C��p�4{J*B1��N���y��IͩA�ī�ta*R[�eF�o� �g����!:ҥ#.V�U@!��3b6J c�W����F�B0D&�18�A[*����g*:5<Y �U�����<��v�ٴQ���w�tG�_����h��ݞ����{�t�,��}��Na�N���c�Œ�k�3���T��Г&��hX�F������x[��aY������R��Ʒ�(FP:?�yZ�(Re�1���̌���tN����Ҹ�2L�nl[�ęt��A�{/.���:���{q#�K���)4�h�7&��� �*�{p����F7Ӻ��H�V�=�h�O����`���r�� �d=��	���a��%�����%`��䮛џ9W?��X<���li�]����}Y��۔$`4P���:Iss�4�I��E+�&�+�J)�o���8",5kKz7Pw����A���a@I���ey� �]ٖ����҆�m����D�g�a�*lO�<^k�@D�A�3ޛ'�Iz�!�k��p�vkӘ�����2V3��Yx���2��Fo��䶀�<�"x�"�t�4�����~��]����^�yDD�^G��.���*�'~9{PO�0�-ӷ��le�aD�P���''�J���3i�D:"5��9@=j���G~��`�� �,D���y�׸��h;�m�̫��v>�2(�&9z�=x����n�(m0��8;-z�v�{��f�O
��iI��B[.ZA1��9�e1���M�2T\����B���.%k@T�Sm�CO�������S�k��[n�eh��A�Ͼ���P��{����R��/`1u����fr��w;�I��Z"�+���p>n#�9~�ڂ�ŝB5��=x�I����G�zA)�Ϋ��6�|��"����a�f�:���P+�����I飉5���x��j0h���gwD�w!���צ�}�ɂ:�w�ɶ2\��n�+��c~/�ħ��ʅ-�n��ƥ8�i���$Nn��ŋ�O3K��Ԏi����#ңI�1mA�?����YM�t���%׷mN�"��SW�W_�,AQI�O0��!�1I�Kƈ���-n��1���Ʌp�Ot��8ƿ��c���c�IP�O(ڲ�Xi�-R�B(�P6�SH����Ѿ��Q�&�"/,u�\�dX>@���d��Gp��A��]�4
����n��dh�w�ͤ���N��,k�'��d*��9Y�t��_4���>��P�xT��.~aB��M��M	4��4Ç� tۏ8=��l<+�����H�4zdS~�h���hp�.�7��'E�;v�.uB��g�|@���N� �� ˯���z�h/"��w�0�x��[�~lC�6k+aц�cH��X���^�q6rZ��T���FM��<U����K}"Un������i�${�h��gs9��:�6�ŉ(��n��qon��͌"i[C:5��41���t�fܷ��So1����lހf��*� ���z��9Ɠ��hũ���S]���SVzD�I�RL�"�yLw�o59b)r�L;3��-ĕ�R�5�6��6����is�����҆�|ZMn��u#w��W�5��u{�H����]3?}�u%?�,*���@��5�(������L��]c�OA蟹�`R��t�͵	���Y�t\��`Y��i4@�E���<�ϋ�w65��#�=���]FЈpH�W����I����cf�����=���t�Ex^���{(�ʫ�u�����yYۯ!?���3�,�M�#:K:���q�w�w���6sF�]T��l�]�O���eD��k����=§�H���N'AK�&Zcq�W�5	*�υ�r�T
�پ�I� ����x�m]�qn���hBm]ֵ��B� 1]�?����J��F�����o������A�J�^���ow��y��s;�0�� �UQ�%�"X����>����o�D����������DR� ��"�	��B��Ґ����x�/8�aN���@>Y)��<BX���˺_�9�n�����&�D,6���5a}�`
��'e�/ؒ�O�D*��X�A@ϻ$�E�������8Q�դh��4@�k��$7r��Qշ���bR�T��wԶV!������u?'��Q��I�>�T
�i��L��UQ���;��Zf�}��x�5�4��7�H�(���u��3WY��g�V����i�bw8V�5���Ɔ��a��<��_�I��C
i_��o�Z��ؓ����c0�]܉Q#�Ħ�}��ܾ��w���5o��[E��8J]*�a�6�BgEB/�!1��v��_tj4lJ�:������*g~��d���:Hx�+����$�����m%������}���u�����-���P�z [��q ��V����6(��k�if�PI�bJ��jo��O����q?��HuJ�EN���a-�����U������5��k��)H#7���u���O�8G�4�+�V�Aqe�3��b��e6�☭2�5#������ Ǧ&�s?�bpX)��x�gur�����?B��B���7F�x���
��g û�Ť��C�>��"3� axuAy�|N��{~C~He���4�Ҟ�g�ь�Z���Q3\#aϞS�L]p`��?�	��'H٥Y�ǎ����9��A����|�o�p�S�@)��8O?��:�\����D���J�੗$����3llJt�l��I�b�%�}H�M��F<�&@���"'M_�"��-�P<7�!0��fb��ı�I�������U0`��$�@��00Y��pwt5	{����l���LtXDyͿ�K~��I���5jH�݆B(4��em�6�,�^�V���O7
�2�3���"q�^�*_�����'�Sw1H>?T�����7�/�#��3�����cfnM����.�k�˓B�s궿�U��	�ZA�������:��k��B�0��ϸ���p��vS�[��`Ly��t�G�H`���4���lK���n܎TJ�a)~�Xvw�֨)�wZsC�kmΨqr��*��K�zl�����m0ę�,�B�-�l���C��W�H�ù��A�pA)LMu�Ћ�b�IXu�¤
u�XI�aP�N�q�%Ԉ�	�O�cK�.#��(b�չ�[�I��JHb�dc����1����dA�a��k��d�i$���Ԥ��7̫7q�D��Gxb#o�H��&7��?[z{o���]y##�6�ߴƩAm������!��H����dg6�ݝH���Ez��0�w�*�g��Zv���J���
�^	�l��v�2R�SQqet�%,�ʫ�h��&�}�yi�ϝu��۠�]4�Ae�e	���AĦ
Y4�t��ے26YK�}��a~��:�~���.��PR�I!<,�vDOZkY%C	L�a�ˬ	~>��E~T����g�Shs�$}�2_��֞N@W�EY��a{#`U G�At�[ �+�<f{�&c1ύP�U�UQ;3g���p�7�`� t�Yo�O�^�����N�*���6�hzDpA�A�	m|,�}�@��6��rzD�s5�����H@�o_U��<(�K�G�He�t����� ���ep���Y]��f>*u{d���YE���O
���9��خ�w|ʀ&F����jzZO ���T�!�*��|{��P�9~� )#.�Uҷ#3}��:%�5�1ݓAI�L���X�j��4j	�*O��� �$�Q÷gw�4����c�e/LL���dw'(KHx�ښ�V�L�xݯ\��­�a����q���Я���D��8���F
Ji�JEzCk0�U��-��Zf;��o�	L��f��|�.����[6��QK���&������b[��+<R�	�ދ����gr;U�P�� ��wUk Y>o�(���V1�ɜC���Q۝��3o�`�3T��P>��� �yg+2�Re�q�Q� �rX��h4�:s[�^:M�=�m>�΅�L�������m�}�z�bڣw+���t���-#)����U=�C��r�It>t@�<~RKγ���Ɵ��t
����B����x<��9P�5�W�6l

����<��{m���%���"�&���U��Y]�E�~�vk�R�>�ƭ@]i\��Z	�c�ēd�ޝ��<MGmcq����_�Z*��he�s��GnR�y��^h�R�Yo��ޫBu�6�R���$��ݡ�9�г�$����*Wu���Ի��.�&ΒJ�ʅY D�薟�� ~N+�znz����S�'�|��_�	�.r�-�F%����(�Y�.�"+�Ó�Q[��O�;�ݮ8�����[ʞs�X���OC���F_�jе٘F�@_(�#)� A~�	��%ve������__��X"��(s%��4\L;��
��(	�+c}]�L�[,E�_�|��4���
���i�G@����}g�"-�oh=�<�sMa?1�'�:>�JP!���i�fm�5D�K3��U�x�������UВ`�?Yb,�W�P�AN4�Z�ޓ��m�MI��*�2��9�Z}�D�#���g��n\�<2ׇ��b�a8�*�
0��؊���$,�۽Ή������+��0���GظlA�ý�����G�V$�'�?(��)֩ W�,}C�lF�]ǻJ޼Հ����( ��@$p�" ��.����j���g�0����Y�7�v��k���,'Z��X�e��/����5 ē�}���$�gN}�3���?��=>��|����	
QS�،S(˘�Y�;phׇ�>���� Z��z�8�I�_t�	�x&q�Q���Iɼ��v�עl�]�L�Q�gD�/��y+��ڔk
i4�2������^x"�x���CQ�����h{�o0���A?h[�\j�ݴ��[�`5��|G���'�i�|C�|ܧ�Y?��*����<)��D|��U� $�	nr*M�*t6SM�bNB?��X��4>� ���r��!�o�˛��>Knsm=��q��R����)���"�4jP�f���<�
��3BXah���4'��5�"l�Ady�\��ĊO��:�*}��;av��j1�Uwe�CE�o�H�e�z�"4(C轍p�ir���_����M�BY@z����L6�0�	���gՕ2�,�L�|g"Tj�~h���s�M�!�х�\=7ts��PI�܅H| �l'�����z��OV��6ڹ�Q��Nve����	Pc�ׁ%�>�.�8T��ʃ[n=r�#0V�����ӹ�v�K	��ǝ*�`v3�����G�RA��"_k��Q��h�!�e
���;��_O��1'i���e�_�i�JH�_��(�a��bVcM�TZ���������:�o�2�$�����'E[lƞ�h	�f<���\v]�`���O���u'�&
��M�/�Oz��I�B
��� V�J�_���QE�ʳ���O��s��k�E��!����*��>X�Ӿ�z�?f�)�Q��C��u��� p�K��b�i#4/�|�.K|o)!&{Ҝ�#��E���KU�R=����`�z���c��N�����Q^���=�O��bM�V�P����C�y�M�@��=[�ê��[B��#���x�'��ay#�A^�����S
e_�9�@�a���o(R�k
L����f	����A��I�
�n�Ob�"pڏl���τ��#�}��k�L���s�t�i���gB�)x���{���ء�F]ϭ�,��J���E��ws`�9f5�"�g�D����� �;@]=d?�����H�a*w�ǘ���,�fQ��̜R��އYP��=�H��3$r�$<5&��_a�O^��Z�P� �4Ϩ��#��j���sj��y�"�H�q	����Sr�¹��a�*:e/�ħ��,E?�w����2����2r!���Ҧr�ɓ9I��P��Rkc�J\��x�+J�����-ˋŸ��`΁�Pg�%��ڜl5��]�j%�����=y�H" �_�Yjz �y:���f�����:o�D$�����o�{��|p��&]�s�H�H�S�j2 �lR���.��bd�l&��}vo<b�@��7���p|���ϟ2��,�9�۝��"����4��5{��q�o���>zB.$��W>&z���W���L.)�H���^����~���͜7u�噬p�o>�)Kɘ��P	E��Te�7n�cU�������N%c�Ϧ�t�i�ғ璎~ϴ
��-�.Ɉ�Y̃H����/U>R���:ӱ��UMP���P �,��ĥ��NU�m[��,է��i��ޢ�s+/3 }ju@1���/G�p�\_��@�ET�Al����bq|Z_�+Cۗk{rߨFr�)��~���3S�2&hP#��$Co���%�Y��D6/�|���0�gζ�>��^d�iR�t���֪ʹ}$v&�`�e?��қp5$as��>��n���-йk���z(F��[���J�^+pr5�j5�r˧%��_�]�=F��g�:J6n��
���/�� �>N�z�{�)
�ama~|��x���3j�$T�\��?Ϩ��	����A�{��W�(���N��$)/�c��;qG�i�Y�k �ul(��|�D����'����\���O��`�X�.����<I$��O	�uF����g�e��u~�_	���lg �Rh�����-_���9��)�	��{O>�Tw�S�W	�ZQ}|!�A[�i��@TfT�R�v
�x��U�n�����K�)
��j������+�����j�2,� ��s�CQ�ǟ/�+S��g�_�T:$��硫}�#�����9�v���>��
w4�}?�@?�=sP�
PN��-:��d�{�Q����s�S J���ۤ�8p���@�r��ټ�X�KBhC<[Q;�)}����;�*�ߒz\�
n���� Yg��N���w�X4lƔ�Y�c��݈@�ٞR��r8	�-������Z� BUO`�u�|�e���K:_�^1e����GX(ӭs�.E��l����Zm�����H�#!3S5��F%Z�iT��!Ŀ������Uazn�qΨW��Rj����'� c2w���U�Ƈqn�Z�������
닩%o $?:��aѷ>�#~�|�C��a<�+K�$?`t�Z�j��Ɩ���Y���A���'7��|4��0�H(��a*��:��+<��,�#�)��������<��/�H�
�*-ʱ͊�K(z_(5��,��.O�jX3��l�e�`�9|���+� :9�--Ĵ���A1i �ƀ!#�3Ũ�3�y`�����\�7'�_P��a��Y�zI|�:�v���`�b��I�׶t�E��{��s�j�y뤒�B��E���2+ߥ�9ls��f;��2p$o1�!\�p��X�z�>{sY��<�j�f����5�4W$o� ��V2����=�Jnb8�!��Q�s~,f\���<�JI��[-H�(�r�Xc�����	��(�^#��B����"�I��n&5�S���������l5���_���"��e���{d۞%�;/@,̘���Hc�C?m�hO��~A��#�.�GW}��^���p����7 ��0��c��!�RP ��!�|�Y�.d1~
��{��~�*�%It�m�_�bM9��3K��<+Kfj��o���,K�oyzୡ�B�����wh�C�![Thl��.K�F)����L���#��q���&�D������5y�E�m����m!o\9l�>&q��Q�t�jԜ\6�ݦ.�P]����B͗�k�^��ݺ��?�7v��	���"0<��V��6��b�ZJ�Ӳ�Z���)�- �-&������P	��~�y`S:�hm�pR?�N�	��v)Sa�m	�N3&Gm)�ge���y9������QE�k�;^��e�wأc�CPM��E�ͳ���l��a ��8��?W9LW�1J���j�\-���S�/$ޢK����~�S��2��5g�ѻ���߂�����o��~Vԍ\�a=��ml��і���C.��:}X �+$[%�W�x�w��3�A�g�C�\Q'��i��y�F05b���ۦ�+q0���wu�yf�r%_X����A�dk�$|�� ��L2j�7��D���
1�ޭ�$�V���	L �e�/;F��OE˓�����Qu!;dmu@�U��,��i��SZ�])�Z%ѥ;%�&�'�H#2����-y�.B�0p�ֆlӭ
��Ȗz�{�)bo9Q��)F�֭���y�H�(ص��F��S�}R�u,�:�@/%��>����d���Ɍ�g�0k;�I4��w�D�a�N�[���]\M����j��'$*o�k_0Ӿ�s撌���Y����|���Ƿ�! av�V��B�h�,L�Rѥ[Lq�A�k��n�RW�'��&N�� W���Ϸ+�K�eD�@+�@�Y�LAd����J*�߇�?��"fZ�Q�i�Kj`�.$��	��Q�u�7��L<}2@�7��4�j� &��/�򝶠�y=\u�����̕+⍼�b�'a� �7�{�I�B���@K���{U��BY>V��Cs}������5Q/:/c��s�Ǥ���:�`�QV"��AAX����U�i��J�j��<��#�g0�ͺ�A�l�ı�؜1�����ULг!�(�")4}nk����T@� ^��;���}�fg��<^Mi��}��y$����8��m�W98J��|���0OBCFSL�|5��,E��8�
R�?5Xvh�~^kz�-L����+Zư�D��Z%"��c�&��KE�tU������Ñ_߂ة$�I�m���s���5��	��L�%�	ÿ�lS��Hf����7�7�2A��`��y|�_W0��rg����X㰢1�e�db���������c�Τ6���7���f|j*��"�P���]����7���`�*)�f�}�Z�6�掤(DQ/V���x�����v{ �p
��d#I;b���Χ���)��xA`|b�U7�
"�\�ξ��#�	�k8U$�ے1��z�>#B�gWu=�^����5:-�i﷞���`4���l�=7�� -�X�㻞����N�)��zU�^87v��B�Y�HA�\<MZ�`�`�8����n��@}�)p7�Eui��s�FL�h@=3��T��VЫO����F�4gA���_Ko�q:,����{z�dof�wY�_ó�3]_����[�'p.��.��m7��h-Z���e�/zf�V'(�������w�ͯޛg���\�@�E�kj�v�K*/<x�	�������s���'�Pw/\��Lgu�R��䬴�Y�7��|��s�m�q��(��F�ٽB������눮�(�g1��k���1��۶u��y0<�G֘�~�1�_~��pc־��ͅ��e�W(/$S0�#�@���%so���f�-���=>%�h#�	l�AbJ��%z].8�< ݦa�mɺ�65�uk�@ �Ȫ��D�I���B�D�Nu[���x�y�JÓ��F��E��U�;��c�E��߬��!)��B��17�ej����{F�������	�x8q!�e����8�e���MF�>�[� �ۈ�c��C���|���bk�CbJoǷ�J�����g >^y>��jÎ�u<.��@������9�Y�ֱ�3����e���p6�L�?�x��@�ɢKל�$��ar��>��0g����˃@�Cv��D�t�e"�i4�V�H*���1��%��0�w�-dI�҂.ʚ�@x>�M/�g����9u�ܕ����X2�.�G`e�=6�����jB�Km�"�=���������u�n0c�!5
��v�1�j��j���;<�Qti7�P���am^�y�����Ͽ�������z��s �Ǭ�S�Yj��B=q���u@Be�s֪���+pFo4%��>�=<HG^�h�J���~d�~��U�F�~�\'<�H���AU��]K
Lmh���n�sM�B0��ʩ${s�����?m7��U�џz&ꍯ>��P� ¡hH=YU�J	t�@����I�X��GOs�F���轳d��ɧ��$a��=��k$m�r0�`��1�f6+���J�tv�r�?�9X����U�'��E�o��JE��~qwcs `?�Q=;�ˣ,*)+_��w;s?���q�ݘ�?O�>�Kj�	 j��^�C�;�^���'��Wr�d�y������|��Ś�N����ְʜ5C��k���Ϯ ��9D�΍���D��˸ʱu��=h���}���7�7���f��o¾��%�&���턹�Y��P�N3���E���,6��lf�[B
�q��N{���g�뚋6��u�`}�h7r�I��gF$4�E��?=*� F���E�0��w���!�<����-����.u1^ʐhquq���X�%����=Q���I�YR�n�s!9�C=�`9=�.]X���y�;>��&/=
&mho@�{���^��9�J|�A�e�;*3,�T镵��!���1���_D6j�4��;&2���>�!;���?�_4��%	�ÈK�Y�̑��(A�|M���EWA�1��T��'Z�kLcp��:ˇ�ɕ	�إҀ��+�wz_*RrɃh���4�I�8�[6����f���}�����]��TL���6�$����M���lfe�D�c��r��ȵ2TW]Xz�Xe82�t���5�f-�Vʘ��A[�+P�^C)����>���:X�Q��h ��	����%��7�sv9n<���� }K6�5+�(�@h��Ѱ\���'W�y/QĤ�0�n�ѫ�Q��B�>)kdnP�����H�W�|���ZN�}��j��Y���?i?"�7HPF�=2[��bڼ���� l}�Y���J�2�s�@2�b��E)A�<NM8��暳ʸ�^��J�Bi��Z�	���+NB�*�����X���?�V�}���ع]q��R d��Y齌���֩�:9fif�TI���QY���g�	�c�G|���#��gg�㳒�ٖO���ω��ŵ�˕FZ4r�L�R��x�h��B�����J�8s����u	�Cf�9	X#��E�R�4�����H�q������C��� w�f�g{N����q^��F�c<#�Y�2/ݬi�� �L 
I��x0/��+M#�f>X��z�50����j�B����E�)�'S�L�[�E�1K��½���*ѷ���(��6|����~�JZ8�2V�ѓ�\�0��6��e���!K�3�%1�Ӊ3��=M���i&A��Ķ"e���t�q�+{�2u�u{�շ{���0B:|�l͘g����;�X`[�\�4����t5�)��A<�;Q� U�Fy�WN䚡�K�@-�8���w͖p���@:ߢ��I�V>Ud+�9����a��rN�Fb��vAn�Qg���X���	^1W�L|r_�]�����@f2D�&�Ale��h&��m��?s7%Kq���x�zY����EܚE�7���P���\e�Z�6�E��eAm��|*�/7vy�<)�et���c��̵��L(,L�٣�@���E���*lo1��u(ي�Nzq���)"�rijDt�o�]��hI��/Hc�ˎ���v�F������90'��	�"BpA3O�q��&wJx]i)�LoO;�ne�Rn��.
%/P���kIL%�$m\؏�2�$Z�b���k ���]��=��\~Z�}�+�S�>��"�D)f^��;^AO]�=�J��W�0-'!\��\R���<h�YO7Of����E��N��WO�u�%�nͰ#p�|�,{�I����[�Ne�PD�	d�r#@S��k�-@p�]��l6��o�Ӹ���>�}��_�&�v���î)vW�����r"�4;�Ɲ��PV�0�p�����
*�'b�!�l����g�`؆N����aUK�R����y�-'�*a�vi�lGx���	���Fͥ��BNF�Q�6e�QE��C��߄�]��Yg���,�?�H��,���H��_��am�>�R��_U������/�.<��h3o�����Ӭ[=߁��]� �W�|.��40�z�[c��\`g�V{��ڏ���4b�P)�^�A�W��E����,A	���̫]��������Z�eqRi���<y�=� s�_��%��3��8�*z ����9k}0b�Q���	�}|J���~���UR��,ʬ��C�]u��ѺHs����$\P��]fy�mSp:�
�k���#Ci��6g��Ş��*�o/(ŕH�Q��Lo�Vh#¥
�]lƧy�qH���*�\��)ʣ�_Xڛ vy� �b���=D䳬�6�047���Kvn�"uyn����#�&H�_� 
R�U�`{-�M���4:�8oj/Xc內�%��*��r	��Mjc{;R-��-��"��[7MKK�#�"V=5ط����.`����R��g�tNn3��D �$wS3���0V�rL�ø�K��ѱ%.9�"�_E-�Ζ�ЬL���E�����CיV���i3���)��{�»a�T�Z���� /�5i9zð����|x�z����v�;)M����ZR�E6�An�s����\��@�9��Ơ�m�ėa�2*�fK�k�K=�w	m1:��ew����Ö�b:7My��j��ɴ@d�q)Lx�,�^���3��P,K`��o �:��H�ӌrV 9�kdYY{����f��g�q���T[�A���nm0���}���?q`8���FW"��קӅKT���v��ɒ`u�0�*��bӗ�v"i���=/��ޛ���	�z�{ğ+�Y�]8���IƷ4o�j�l�Φ�K���
��R���٥�:
Ǿƙ֠r�(�i����ma����k|�mxr�#ܵj�Q��
9��8�s2�b3S$Փ�2�
K�y��c�Ҕ�Z�=
��8�+�a�_Q
���i6l_��cndq�����%�� ߸�>U���`��m��Sף�=T��^ rd���|8�I�Ļ�S�ݍ��G�Yʾ�7�:f����6�4���jʽo3P�����`5z%c�0$�o%���%�}�T�8K�A��\�6�n�]�^ΞZq���<ڊ�l�s�+~P3��rU�v&�L��qX\�\|���A����E��u��g�E
6��V/�p��J���&���nn]��E<	�x����'k3�>;��ec��L��ݪ[����p�Kvʹ=�vK;�����z���T��fa�n�_��p
ۏ�����]	sT��쾟���g�zJ!�^�et�Ic�@�g��c:b����
��w^���}��h7}�h$`�!j��W��1�t���u��$�p*N���X�<�n�B�P@CC�(ߐ�W6Lb'�h�*�{o� �?�@\��c
 9���@�ɞ]�%���� ].�i���C侎�kf�����^���+���U
9�G�q$ݺ��-B>�(���=��ƕvť���#�(5�b%��gK������zSA��Z5���';ӓHAvI׏�M�Nuy!>�pQ�B��u�_8���c@�����"ӭ7��聃��$BC��ژ`0�F�hf��67�b��wL�.�0�@�I���j<�?��SZ�/��$|N�1�����չTt��ʥ��;��]\a��g��kU̠��I���g��_�z��p�t$.۳1��XFOT�#P+9��w���B)��B��D�(���T�����9�zS�Z��é7u�}.pn�m�4}��G�v[�Z^���;���[P*o�����z�QC����Ծc�w��vT_#Po2��ʪ� �݋1��*�:���Q j�4��} ��0Р�(�OCd�}6vN��Y:GE��>�MJ��F������N��d����T�߅�JO���`��F�Ήr����f
+яhN��d��y�t@�p���Z�_34>���B�q~�bōr�0�V��O_�χ��C;�����-&W�����������S���<��gq�?�˰u��9��H�4۟%���ٺs)�D4���v-�u�Ǽ�1�{ Ff�o5W�&��W���p0��4�gh'$s����MS�l,�T�3�M�rl?�_���="'1���ثh(<��o��z�){��i:�|,��-)o��i�v�� C�GK�J���`Jh�K�X��%[L1���q��}<���X�)��CT�o�a@���N��^;��(�9�Z���:0]0�jC�X�\1$\f�N| "�&�X��H14�Su�����#wls���*��x ՜�p6�|�����$,_miΣ���[ھ9	��-;_{8�6�$,�k�����/�m�{[w��z�R �E�tK>qR�6�v�	�g�L�_�����>HQ{���"�%Z�FM�j
�� �7��ٞN�:�uQM��4
 yf���֏��Z\Bp��`ih�Z�΋��s����_�3��2�ޠ����r��/�¹�N��G=�"�!ć5r�N5���Vt^B8������;��e�X�FI��A'���T�gߘ=Z�ĘN��� �(##�Or��q��g:�>��ԓcL9[A9���㰄����ו���<� ���v�5�#[���$ap��~�,��'�_���.K@�'��z9���uCB[�g��M�L�/A��H���8uw�ިJ����o:	�4�e�P{�3`�,	'w�%>����ԫE��Ǉ��&���Z�nIȥ6$8� ��}H?�3H�0p`2'���B����e��(�I�P�cay���'��������v�fp\;|��Ȱ��5����=7>Ȭ}�r��!�ب"�ĝ���3���E�Ai\>�s����Ĝ�3j9�K��m4T,��ϴ=9����pXQ�$Kh�A}���js�ު��b,���ЯW��5'��}��i�w^��g�Õ��Y7��cn躾W;�${�{�V��1!�Ԁ��k�	�_�����J�}���P̋[STl��O#uu��C�4���%�k�!e�D�8`y�*�6 &��\�!ާ�9(�'p(e��+�y�K`��ȅd���0��K�?�n�i��(��ʒ�*Ob����S-Ne����R���g&9��"�nE<4wC��Zũ�L'>|/3Y��5z0H�|X��Pu^*�g��#|�^��Q#��n8S<Q�y����$�7pgFE����-�p&]U��g~ �)<� ɗ�������Ֆ{_6.��ۭ�C�L����+6���N׭ƽ����paZ|x!Y������|�5�X�q��/�bz�c���D1��}��� bc��G&܉rg��7�۫_�
�u�&�"
E���|�Z���[b�&<p.B�i}�3�e�vh*��`\T��0���w�i��]���U⠇uN*e:k*��:4O-2��4�Uu�ˊ9�;���@1h%c�j�6٣D��/�_�3�,2���{��?^n]4���O�(�-7�}�}<�ü���Ks_��Ů��!�J���bB��{(&��¶�����I����@iouqs\���.C__�]���|����?k�؊��Y4^�d����w��)���QY�������B��F]`�S|��35�A�Y��	�-����3��=+u���/��ไ#9��~b�j�	�I�O[���q_/�t��9�?���=
 �'ϟa��5�v.>��cl/�f>���U��1/�o,wr��!n'����p#��N���ي����e�g'Xa}�}��mz��
���x�VH�Ǜ��f[��Oy*t�U��i.ۭ����ķ��L%��z�bw$��N8A%�j�&��nF|�~��w��<c~���<��DIS��_�& b]4�b����/����l-2�������H���/f�<��ѽ�-���&Q����&������U0���Km�.�������^��^U��x?���b72B`�)�Ab^G��4��ȧ��L��9:�j�����?v�U�<���ʯ�#u�7�P��u��FZ��
׳j���۳��#��Gc	���5�䖰ݾA2�V��������ٽ]��|ۛ��Yc��@#M:nFáa�]����fS�������?ڳ�?�d��5�$ꎟQ~�uXpU?8(U. �����9�q^�kl=|�����A�d�b��S�z�2Ν��ܾ7��"�N`e��(i���!�Q��a��4
OP�;��J��R����i�9�{��2bF������J0+Vӿ��U�4t���jS}_̥A$�Y�6m��.�MHh5�)�+!��1q��ۡ��=#?&����M��Ul	����^�ɭᫎ�z����bu��K��Oy^�+s%N���	%�$���FrUa<.+�o{E��zR�K>k�ڐ��Tl~p��UF^5q����$܆	#浰���T/>�GjHE��M#������ܪ�D<u4�o�b�ʑ�������d���iV�'X�=�OȬ��!?=�E����R����{��n��������T'�ߞ
���#�/��WX琧���y~;:;�K�5^��gW��bSf:� <�LnJTe�r��X�Q�A������#�ͩ�5v��,�R���K��ő;�.N���%C�fD��q"�]fV�䇤t&>~��Y<�6��7�gB
�`��3u�	Pr>7���`fu�ִ��y�)A^��՜1P��|��&:^��NM2?����6�)	\�Y���8�~��[5xi�P�s���{Ѳ��K�;���m�%ـ�][=�*�9�(�[w؋��.� 'Z6�F�f�`�����}����`_�2W�Z�#� ��O?.�EAH9��H�1���(X�x��vo!<���V�sJ;d�]�	N�Fhb�C�+�B�� �c>��.�c�;��� ��?�=���%%n*�C��מqLUu���+���b�f�c�Ǚx$���`�}���V%$l��8$�"�#p�|�ʹ�I(���Vx��jn�cp=T���ψ�@،�?�f�e��B�I��p&��'3��,&	9�����#���,,�����D��
ln1�,�9X��D���_wnTx��ս���T74*��K���è��b.�DV��oF�S?��4O�)RP�6���Gx���$9maJ��&��㡭i=��b	1� �H,F� ���L&-���g�HOW"�q}�pR����e�795�G!����+x_��8�2}�]�#��Ъ?DN�W!�<��5��:*�K_~�l�i��I*�ʫ-�y���)�����ۗ�n�[+vӯ��R��~�U�$�XJ ��\��)vO���;��MT�dE�s�$>��1?<�����p����0�╇��Y��^<�mt5�jo0r��w^�=���n����vV��8����,�hz�?1�d5>˂�����T�L[Q`�V�/��<hOmph$i����:f�)���K�=Yqb��Ŗ���UY}��t9khۡ�a"���v?k|�L����׆A�kOŐɌ%���p��ƶ���5�pT1��c���^��NP^$��	|�#}ϗY�-�+��vu�ij��>���'6����D&��Us \�E��� �y��|�u��wH��4�i�c��4S��n�y!����HI�������~���C�f��ፂ�o�1En�/��={�P3󍑶��Bk�U͚�i�;E��
�G� �S"�]U{�q�ѭ�g&^�?`��F����ǹ�K&����Ն�'֚��S9�Ǧ+N���s��x�F2>&y�D�6�LE�u�� �3D�OH?�ٕ�j.� 8�y�s���\��cB�
C$[p�<�{�u_���9�F��0��ӓ�[�A/�sI,��H�`\��|y1���D2� Ă�CL�$޵KJ�w-�V�GӖ�����=E e�Ib:.�PC����8���E�̷̩i7P�����k�dozћU+�����H �M�G�f+#��4d����u����g�O���0�	�y���DJ�-�vl4�Yͭ���D�) %�z�1%�·&D�;,P��˿��<�czw�WATxh�]���{v�N�Tj^��_��%a�9�]@g�6�����b�3So*��-Q��f9�n���O��}��W䜅/]����m������Vא��d�k?����6%����AɢV�ʠ�jKq_}Ī��lKTi��!�S#�'�q�Z�xl�p��&�iN�t�z}�@61��yR�e�B}M�}j����[�0��.	b�Kn���J[�hޡJEH�ldhߧ��ߖ�'ˀ�6Yb�F�K%�w(6B@q3 �$���ʈ5��E�B�s�Ԝ+�a�6��İ"S f,�4)c�)^1E�iMގٓ!sF���q�X��o��gM��U�:A��IJ�	تu�|�����l���kWm��2h�n��s�����Q|3��{��x^�~����m�R_�>�vE��w�ח�զg����K䘩�'��auf�7Q���KS�ZG�]�մ]�5��X�֓vm���2zлG3{��[�($5�f)*ZӞ�4���ҧ� -8N�1d�h�B�
�j�R��.j䅌x���,�9�5��aWD.p$����>�m�qSH��'�R+�]^�$�!Z�*e6�7��->��@V�|SNv���G�ݖjYҹV7j;{�rd
0�bs���)P,K�f�0C�9�?�@�>_�%jU��R6A���$�����$���� ,l,R�y]����oJݣ*�U/qC�4��)b�Kd�"k���*`�b�	�9��H/�"����ث�w��!�:5]�#lL���9���qY4�G%�VŦ��v��u��[��D�O�vCn��=;97f��KlGiⓒ��"�>R8�����pv1�
�����RPd�,a�<'�0�����s�w��k���J$���u@&H�@����H� �P�쑍�܂�l
~Z�@�5��� 3���D�'E�|U�����6~c�ߔ���Ň���0�[E}���Br��!s}`���ͻ���@���|m�q�UTI���7��m/;0L���p�g��T��ڗ��Ư����?�{�d�
����Cu�/�X�=-(kT��;E�s����TƴϹ��UšS_�yO
6��p!#d������	�Ãn���+�FC)�QD�16�)w���2?b(́�7J��ż�h�{�8�y@+U�I�ތ+�x�����.D�G ��
0���D[�NX'�uh�#����vt�	�<�>A�����}��=�~u*�Q*�r������|];£o��//.tܞ��%���w��;��p����>��r�,�� X��&�׃�G��zDfĪ�%)�)0����	�,f���s�)��ֲ�IN�C��'�`#�c�%'�Gh��6+�����s#��Z��A��D�yfQ����}#�aZ�����lI6o��2��_�O�s��P���Un}E�,��Ԝ]�}V��h�)�!�RV�M{O��%`�$�*�?or��1�〫���7bSα> �i����Ce�l�v� ��t���BR��_���w�!�������Iҗ��_&�|�*y�U,D��M����� �,+,Z<	{=d�,u�r���@�)�l�G��r��P#����6��A'i����ٹS�<c��|�8��"��T���N��S��1�m�e �Z�w˼e����\BF�C �:��v��m���p�0��Pv���F�ۮ���9N@O��z�����y���ƪ��@U�ʘ^+a��9���	��X8~��y6����������V����ؘ蝓�8���RWz������ ��i5<�2����^�5Dp/������k�� t�L���z_)�I�y˶��sT����Y�t�_�J�,'2����N:8&��f�����᱁d�`��ʐ��R�m&�e D��#;T�"��<�>W���8
g���(�������H���!���v*�;�	B����y���K���Q��i.gI͑S�-j�P�c�k7�?w]�a��F|�!���dg��.(�͊�}d����$$׬�t=
��Z�P�9���# a�T�s��w�Éh���5n�D��ۨ	�:�&v�*�}�3�p�u��)����7~���Mw]ɮojٔ��v�z�`~:$����+��2S��:ν�eR'o��r�׈;�w���^�~祳 ���ZSn_l߹�|r��"t���|cp��g� I$g)k�#j��>�~W�_�+IlvJ�"I�ҫF���U��#�Ab\:�'�h6n��qO]��Y/���3n��膶Zƚ�E\�P��NL�������8����|7&c�WH(�P����Ϯ�	��E�A}NKm�A���}�E��?p2J�SҰ(ԯ,��:�L�Ĺ�Ű��34ω�U���>c���#x&\�E���@�!���@�L_��Ax""�΂�z"^��zgXY���N$7����ċV��XLN�.�(�Isqr�8bFX��#��}�^�8��ۍ�Ie��?��S�`�^[3�2��h�_���)(��]��L�N�Ex��%k��}x�z��zT��צ�{�<��:�L�����͞*�F���X�DF�c#8��������:�����k����elГk��X���.���^�<6x7�R;U�Ih��Vqؑ,��D���(��U�� a�P.L-�(�s3��%_���Q�ѻ�[��Y�� �"'�{�VFUS4�P��~���EKbgZ����k�,]���)gs]��
G�K!�%�4#T��T����q���OI�(R��[����!����N���^Z�Zd_JKXA��$�un�p1!`>�>�y	������I��˃��c��ת��&G�@�5L`�a hD�)�p��[[��^a�(%�/V�T�=��],!v�J�&�E��N�ցN�_�$ă��BD!V����\9΃��3���v��v�'�ߘ(�Y�*T���qO_~��S���<�Fܛy���Fn�Bve��fs0z
�t�0�Rv�^h�i��"]߸����y)+li(���fc��M�ɩG�Q"}���X�\�O�QB��Gb����}��,\]�XGc�wUF������њ��n��7�J�3(89jiҎK�]z�Qu��L�S ��q7��W}3�YW�ݟ�?b����"�K�]�Ɍ�h(�����u����Å<��Z8�k�ըH�&�+9�X�pAO����`;����nG��E� �BeX��)��a�yi���e,�	l��8.j���(�U�ƀ���h�J93ޭ�FG[�
Sqb��������z��Dx[�mXe�a�>�:ӄ��˦�jc�k$�ֈ��~0) >�h��ư@��i��|t�4-�x�v���6#�9��T|o�3*�G��c�x�-�3/r=>�A0���w�9�W�Q�����*/�A��>x@�[��^߫iևݐD@��jȔ�}Tl)��3z���~f+���9�o����_��yR�J�s|�~��b���:"�������[+�`�eP���T�iPb���R��?{xq�"i�+�����4t{ #�7�}�����x�c-��w�
����t癙3����ʭ����
��L�̭;QZh���0�(�y�21�]��?��W����Me��kך�=��$b��%�1c���Qw��b_!����(��������l��eZQW@S �v$��kq_B~��L���P���z���[۲������(voS�1ᴸ��_b4��f�v��IY�na��&���j̻�N��J�����2fy�w��q��VZD�K̒L�DDض����\c�����A��:�D��F՚�O˞sBo�I�U�b�S˴��,�����L�=���ERHT�#��@kN�c%������O���w#Q�`�B�>S[9p!H��?Du���D��ֿ�9Qyqş�����֧�Ui�A0xh]���3:gE�*yXM�? �$?��rF����:X����(Z��0��~��>�N;��y��Q-ڄ|�^�4�M7�/��j4��3)b�:��-�aG`>�Ә=G����X�JJ�p��X1+q�|��F����Q��
���)v�emM��pTێm2��!�3�ն�����)"��<��)�����D���KTC���ʽJ2�d���ȸf�8w��1��qźc%G�B�'���^� p�y^W9z^Iڅų��m�0��"�2��dƜS�I:� .2���B�?i^Ύuߖ@3��ƍ�<ӂ��'����7\��WN��@X;��	�:z�F��KZf4�fn�
�3�	 k�����l���>�u�h-����t�;/\&۵�X�^*|-�L��F����b3P#l���6�W�=/�<�@��T5����g.oy�Ty�o�P^�}4��Lo�M+�b=x�\2'�Fc�<҄k$�"���0f�GH$}q]����^�4;$
,����ru�R3}ЕV�dN�+IE��ؚ��>g�F��n����2�� %���H��S45s��TFzB_�~������{�Ly�,�@�&>�]��"婞2G�Q��7)����@l_�վ�T
�KL��4(tȽ�c�;sk���8���n�8|��"��U���F#<X�V�1�j̶�1
Ί�ox$��D�.U#m�4�8�@�/��n�!)�sx�U���$o4q�5���@1>v����vI��� �m#a	��4����_,��
E�ձ��<��L�:o��� ��{ ��Y��/�����/c��<���	F�]][�[��.�;m?Ԣ.`bLB��s���攙w�����;�m��+8,ټZZ�_���C���Ǳ6��Y�������/e�};{��dY,� 4qu�lr�$K&R�:%��	�ׄV$FLZ����,�&�n|��"�䢞�i�To��w{���
��V�پ��]	�3�ap�@%�NN5-6C���J�l�Li0��Zc(L���0�0�&��{ܡ/�-p����M��l:W?�z�@T?Tu�,����c�_�gQ=E���Vރ\�h�D�A� ��'z��t��X�M3BTv����w�3�k�HO�7�`���vd�w���|��1 ��Y0�gv�kP���E�IG���j��ˏ��[ӸR���nv������T�@q�VMء��u �k�=��?3�����	 �Ȓ�j4�U����P��,}!I�9i`�u"{��R�hU��I�$`-"m[P3�:-ji�x����=�W�1�w�~�A��T�{�T�n
d%׌�,��L���ݑ�i�n'��ީ��uvgvr���^���y	�&$��+/��/�Ȁ�5z.9`�:־Шq�1���`K����j#i,=�WT�#9���Y��A�*��a=�1���2���m�؞�g�K�UU���}YI���g����	>��/���#]{�R|�bC���Z�j�>��;\���Bcs����qO�W��H���T�(\��I'B�4�/MX�c/���~"�
u�	n��1ݞ�����,g�6��O\���:Y�C��Ac��ӓ�l�j�Ŭ5ߠ��^��{��Z��a��˝��MW����ܣ�L�_�O�R^�[�{�.�z�Fd!����	ڈ�:'a�Z�@}M8����48%���� LEb�Dx�4��B"|hȡ��+Fe^:&Ѫ�1��;;.�d�Y���\�
>G��M�?�V�Y�I{�q����[SO�ý�;�(�m��2x�"�(~&�N�LYF��V.`Bh)5���=aJV~BK�C���<YI%��8�Ƶ��*�	?�����Dq�1����]��e�Q�:�N�1��il�Kآ�Q��U�����Ѯ|?zo�c�R bY��I���o�V�q"}�4���G�����lq�ВwV�A���#��5C������}���
j���w����0��@�i-�C�w/�x@NƑv���M��N����H;y�N��X:'�����d;e�+I�/�P�-}�P�B*M�z2Wz�c�<���>K��>���|�$w��P��qlһ=�1����'�ʂ�FT`���g��2u� ��=�ӎFi���B�d�ݵ1���o�"�s���c�u���.ʂcj�y��^�C�N���((�v�^���e%�tD����� �;�K�^e�7�ؼ̥z��{�$�>f��]s�̀'S����I��ɿ���,�l��U��{���L��&�m�=�+�!�F!k�����)����x����T�4�  &~0���EV��E�_��͇�X������]:Xd���W"���������5�l�ė�F����3�W��03]/���@�O|��I#k���`����&��q<�z�]��<�'k������P�wCY�]�k�����]c�v�h	�:A� ��\_�H`�iH���޶�>����@�D���o����d�����rR�qv/��Ae�Q2�":�ɬʑ'�{&Ǟ�e]��+(�c�,vn"2uh3����5o	�3��>mrn� �m���n��<��b���t��[O�n3��Ԁ�M��R-f��Ȫ��h*y���[{i 70�_��2]�7#B���*���	Z��۶/[���MG�����-�#H$L�5�zo$K2�蚍}��O#<tH�	վ[0�{^ϛq�y�U�E�i%�}���\��F��jeϕΣj���ܯOR��F�?��6gG��3�@���%�����OC��g�:��Qx{hDo�_7���w:� ���
6ܻrK	.=��h�6���8w��G�
�D����n&.om[�"�g����7 )�Ji[� d.E�PE�@�9���+�/3-M<ɘ�>jn�߄sP�͡�Ts\}�8Ni6��5�v�_�� ��6�~��y
 -��rl�a�R.��9r&z�h>����ٲV��� ��Mx.oA����
ASQ��|!��+�)���T���b��;�(�f��h'2Xr���ĭ�jӒ�W~%K�������	�Slq���E�q1��� ���@��oN0̀�<[����~k�J�PH�m�g�ғJ	����7$���R�kz��Bd��8,/e��wT����ޭ��Y��\�jQ+��Ko7Po({���7�N^f��蘼��M}F�|!Q����%�.�X�!�v�&�],2����uS��~vnۿ�dȸ|i��v"뷞n˖�6<��4�E��Xv9\|w.3��@>�d9��2xd1/��Ғ�U?��~3L�-��_OpC�Y�wk" ��T�������J`Uyi�N4��48�K��]}E��Ň�܏<cY�:c']/����
&�$�(�&O�p�ϥ�P����5����[�b�K, a�p������Jê�vso�a³c��j ��I ��!�����w���b�꿉/���S	0'83��	�0��a�i]O�.;Ӏ�9n�#=!�"�)��`���{�|ed����#T��(����=�Q��y�b��2�����iɭF�*n��(��K�ln���m�����r�	���]$�h
 
��0�}�Gu�����!e!|��+�~s2ѠI�I�+pn��N�@ow�#k��L�w�E���?���޽R�@$'���ざ�OCAޱY�}儸�H{��'
�[�0f�q<Ϟ1('�&��� �,����]��s�$2_�c��aDVq���;&�y>�^{���j����������R��!a��]���	,a"�ٌ��(�+�[W�Δ�b���*-5�z�We˫��zE�.��|ٸ��l���-�]�ˬD���O8��]ս�oe���^,�1Қ�(�2M���A_�5�&��=^���}**���ۏ�o�Ih��o�*��]ݻ���^��Щ'd�L9�i-BI��p�V`RW��A���/��s}ͱDM��?��2��' 6�)�����L�K���D:�c�Ej��G��}���_�w8 ŷ�J�l40������s��Y���C^#�j!��;W�I���KW=y,��{D��i�o���ɍ�1�f�?g�1z�~V\�Eƨ*�>ug(Y�˓V�Oq>�,�W,,>�g���X� 4 2���s�ò[`HȽ��7�Q4����7df�7��PN�'�G��F�i^���Ɗڜ#�zoN񗼈��'[B�����.��'' OC���EC �W��np��st�����7
�}^�c��5��n�5���b�Q4}��#R��J8\��,c{"�#ALj���K�k�5!8�Wc��B:,�o�0@�t(\�t�̫��	��QJ`����l����'��w��XĎs��+
V�C�g�=�H"��t5QH���o���>/ࡓ:P�~��==� >Ņfd��Uz��I	f_�2\��r�bo�ڸ��Їb�NR(U3�?��	� � ���ݺ���x����:���2��.4G�ʋ�v��b
K�n�b6��ȵ���%ٟM|�W���ʑf
���q*�^{迻&-!;�H�D
	�p��S��B�P�o�fk�}�^cֺ�"-����_A�7]l�9i�R��y�Lr�QS[�It� ��_�b�`�[Ū�cbw��V��6m.��$�&�I�~)I��{��>S�[)(��ؗEt��E�Փ��34f�ڴ&#?��2V	t�f9ma�:���$�4=;�k�'*�	79���GM�s['%��E��G�k��Wd 	�d��~�Jo��J��]Z_�����m��Y�:�W��޻6Y~�Php�'���ξwN9k^�:����nu���!�1�"O���\Z����۱�ƈ��zJ�m/}#W�x#}��T���R#�̫7��`]X�V�~�G�^߬��;�����v��s'��2�[ԷS�\��4�	��"ޣI��`bWu;�{ĭ��M���K�Ex���S%0.��Ėd���ю�iSH���(����@��g�	!���X�q�h7*63�i�����4w����ϐ&r��[�q?}�	��k���;�:O�,�
lb�ʆs�O���{��04�e*�:�A48j��q�K��̒�L2{d���b���'AС��ʢ��S��)�h����|ζyJ�ی
��gφ��O8tE�砛X�/:�����-q�S5?�����"^ ����f��q/�\~�C���==t6��Q�Q4�r$���TS���3(~�e�:=�r���}dF+]~pP�)��Ab�X�h�g�%yu�(���l,������&F��d)Y,u��|I��O�8H��V"Q&�Y+dI��ŧ0.!�q�԰�"k���֚����b���	������a�� xQ��\�
�Q��G�T��V�,�,U=ʿxp��n��{�LP���*�Z:��������9�j_��%����I2�M#0'�(m22�Dj��W��=Ĺq�r�G��������.Vle�qn���]�Q�L��i~��F��]�LŨ�i]����U/KrlD�2�a�s��`X���CΊ�\ħ�qb�����lܪ�u�7o�P�,��B�%U�J麏�	�Y�$���[��:�y	]��ɻS�SY�B*�{x�ʹrv�s�7fd#�����ؼ֙[M"!��콋�&�@r�#5zx#�Q�un��pf7�s���鷊xu�Y�'dR���[�*N.�
w>�!"�$�O�#a`�N�c�[���A�u�l��B�(	��L�9ˮJe@���FP9���;�EԾ;��c0�Ϣ�D�����9����svC�]m|�G����% 2\�d���A"�Hω"�����a�f%�x fp"�k�}55��@ch�*��Ǔ�xk4nY!K�2�c�t���k%(W��Tu(���#t�[S*��(^>^��b���=�X�+b������d��"�8	��mZ
Ǟ1�;����������$��G9�hQ�ٶ���j7�W����-�-."�T�{J���Bm�"�Չ�(o�G��3l'�R�e����S����p��&iา���I�˱�QC/��;��x�uڭ�鮞�Q��h'E�c
_#:\�BK���`*��t�{�y�Z�$���Q 'doЬ����BZP��y��CV�<�*��T�&>�)B�����-�R��v�t���d�Hc�Z��꫌
�[̸�c�ű��fbE��/�����X�I���OG4:�h��{KS|����Zd���
r��.��0��~��"� m���.���J��yiG�{�C�RO�g��Gk�2���xn�:>�m��̵ٮ:�ow,a�+����D���@���d��O��
�|�w8"�@�*By:�P,�ų1Ǡ��\d�O��+\�*i+��(��(�K��������@IZJ?}@��}���+�-D���ӛ��Kn�R�4�p�'�in���X$�`�����=j��u������KyqXE�_���/p��+����m7�~��Q�X��R�v���J̕č��N�g4дD�\��|�BcB궬֚�Epq�w�_�Ap"�7��0d���f@��i�������
�g2�w���[�U�����/D"��pA
�D��x�!Q����mx����+g/������� ���ve�ͪt4��=0)����h��>�*��Jk��˓,�DD���@h�E)N��P}I���2i7Q6� �;/1��Z4N�����[B�F�=q���'�kIS�`X���ƻd+�COE����h�] �k"{xz*@��a =e;&������������&��Y0Ny��w�T#�c��3P�s�+�GM�ĺ_х�Hg�Ⴚydw�#^��G��Э���i�_�i�P���L�p�����+,�fĥ"��_do"�c�R��u'[����NPV���r���F�1����Q�V��K &�����ip~�z�N�G���]l�K���8Xhfˊ�m8���c"}OҴ`2���e%�Hto[�0`c��<��N	�Cù�}D�Ûp��hg���;�n#@��+D��XZe�k�R�?��P�q�L�u?5�`�9'�4�3��7��l�"@�" ��ׅ��4 �N��Ђ��bk�{�I�SɁU�7�k˧}gpM-u(�-������V!�)B��Em'm�i���E ��.��(��	��c���D������P��g�����
WC����q�)��� ���!;?Rn}�v��=�{�;�p�[��0<�)��ՑJ%x\jP8�f����]G9�'V6�Դ<��5�#)-�
����@)@�Y�a!P��A��𴷐�����,ɒߍY�z� Q�=`�~�G`�
�����vJh�0,R-%�Ȯ�L	wxݘ��"�e H��R�U��&��R@XR���5\E),��E���#���5�_g�E-BfU!iX��xx��ˡV;t�f]D�/�B�fZ8���X�?�?���R��}eN4.2���O)��B��	��u	�@/dӝ�R��x���Z��{�q���X���ѫC�ڨ~&�^�hkkt�.����{ZjX/��g���:1��7�7�q�7��1�E��y�Hyǅ�g7��s�v�P 2
};ۀ��>R����--�yꊅ���O�l����M�4��M����9�j���z��;!�;�0$k3(AN���<�A������e�OIɆԲ�R��=��(�c_���zd�Q�<�Ew��ta(��"_����l������&��C1����W	vI���yٻ0QQ��z��-� t�e��\U�GzF X��k������<q��nP3VL��J�0���+����O���\�N���ɇ`�FcN݄���Z�sQ�k�D�:��<�ġ1d�#���HG���Z(2=��,?i�wD���V`/H7�v�-i.�B�n�����I D����5O@n�ry
a����Iɐ��&RÅ
������x�����Y@�Z�sS@R���(�c�^,��J��hm�e�z��Ś���l���_*�tJ��( 	�H[�fw�I�%�8:�$<0Eŷ�"à��6=��  "�]z�s�<bw,�O�Q��ܠ}�]{��U��o:#y.;�腅�a��z
s@op��H����!��}Q�\�
�Ä����~��'bם.��K��+��@����{����=�lҒB�q2\_T����=և��J�b@�i}��,:�����J�d`�{�9��g������<1�*��t���S	Ȭ�T�D;�DF�;���	?(ּ�h��Hm�;�jCgx��t���3���D\������(tF�x�� �U�g`�=���
�P��iBڰ"�G%�y�����QG��
�ڌ�e&��y�"}L:��y��e��k���$y��/�3x�<�J�W(N+)������-����/֩�5�Ŀk���	�%N���h��{^�C�;�:V~�Su���o��)���Tب�?��8g"��	�$,��]�v,	T	+���E̒�#j�~��g�~�/iZ��s�N�q[�#2��c[����"��q�o� 5J���s����j���a��Z�=���o����}(*n����]e�t|�ӫX�-8-T���'e1��ɥ_�v��h��^oC��3�ג��D��#d�I�����M�ߵ;��'�5Y>��K����o�X��{Y��P�|�l�>�fc+&o$0�@��蕻�5��a~|T/�u�ރ0B�����s�E�۶�46b��N�f����;N��J��) �s��*,2J��O�ku2�̉�)ޔ�Y�]�$�Mmb���pQ�ʟsf�A$�wH���0W��ӭy��<=bײ��\"�!i��H��n����[���l�J�����D  `e���Zu�Os���ES��z�NJ��!����,�ֆ~@����m�d�O>����R{N?��ڟL��@J�#�n5�6�yL�͙�3J��� �|�V��Y��i�!F.O��ݟ�R�~J�M�3��|��l�_1����):�U��Y�!�Bd��6n�|90{ӻ��`|�i�1A�M�
����@�m�JӉ)g �C�Y�j��J".\�j��_�%�W	L��v�	g�����|�zΦ Z���u/P �����+��������P��d8�~*�S���;�*#m�PD9�x�.�d�(*�W��H�M0�Dt{Xt7/�9ڍez��&<T�9�B�N�4b��|�}���g�[�ŧ�\\z�T��n�3�!o��+�>�p'�7��cC᠅o�*�N�v�H�D�x�І�JU����9��OU �d1W=HHk*�E�����kG	aN�^V��LW�S`�4LW���e��ޘ�jǦ��0���(|��r�%�Na(2��4�s�f�w�U�� 8ܠ�m��j
J�.Be�eꇲg�K9\�	��]����{�Q�#[��	�,�._ �K6?�y�,���d2:f���Ko�Gx'��٪��a��di m��ݴ��o$�?�h{�X7�a`3�;ؚ����������k!_�s0��Կ�O����d�Oĉ�Տsړ\����)���&R���q�zw*��K}�q+��+Ǝ5�!x7�|'�[B���y����cR�U-�	%�d�R#{CԾ�:g�r�%�U=��uvN��_~D^&��[V�ʺ�A]�?@E�G��Ƈ����̋mgqF)������6/��7��𳽦#�_o���-��B���a�%�ʁ�{&�,��_�|�:->�aS^�@��0����"V�����qѪ����]���7�ΓJ�^9��R�����-۸����<�DU�~ZzS����9T���!X�~o�<�p$��
��y�$��9z�)_e`
�+v�K��\���f-���ֻ���9�L����z��g�¼-�%fy����;{�S���!��7'���	(�Kv�eެ�@��C�'9PB ��?y�pC{�E��Q+�k[�s��K��R��iH�"ĺ;����X}f�h��%����[���yTAF��{J� ߀�@��c����9�j[�?�,?6��f\i��ajrz+�QGn�p�n�	�)iƮ�BOl��p�w}Ee߳��m
�A@r��e$������0TU��L���H�4��U��M������cy����������0w�����w,*����\ۙ��:�ݘd�j��p���N�8X��Do�a�e��w2�9�!��t��CS�g7T�:B�J���Z�C��q)��̌\�)�y�dd��ӴuȒօM�*��B���U��X�}���րw�i��{�4��[f{2�� %ƾ�Ȭe���#K�6I���Pɨ�ҭi�m��r%S�è&U�)��f�4�*X�D��A%�x�&".��u�=?��arvRЌ%[��\M��9M$<��"��Dt1�xTQw`�X����^+!�7%�<�P�1s|S��N�F�g�.�U���W��L��(�Ⱦ�}5ejuY�̛,80���䋿Վ���x�����:�XdXP��MA�r _`	S̴�.0Y�d�Gݩ��[������/��'�q�

�� �ȷ�N�V�|�͢ߋ�/�MhO��&bl���&��sc�p���}EO�'<8�+<{�[᳉+	���؋���J���d��-��A�i.�3pdY5A`
�&G�Ū��%�&�0:vH}�&��4̟4a�o�*�[W�6q�a,�O���l����S�o����Å^a��U�8g����ȅ.�z�~�
�ؔ�[aj4n��31�d3�GG��wR'zǶiM��`������;�SȌ��
j
}�/�+�bə�J�M̤���Z�{i5�ѡe7~n:��K�+�gf�t�Ǘ����`��a)5`��;bX��J�m�~�U��~z���,�0#E����!����'��\���{�&K Y�=���LD�s#t5�A����s�a=y9��RGVt�lT\�0F�آ=��k�{ݙ����>C�,O�r��סr:�KK#���m����р߿�9	���4���tCI�|�-&�k姬���k͡c��6l��p�K�|����������Zz�S�C%n���f��g�2�[ѐ�����Cۿ��Ļ"�6|E�B�5�W�1�'L��=� -k�K�bϫ�nmK�k/B�c���`# ��g�Tւ����7�/e��MTn��m�d��g���gMs	q�g�.�CQÜ@T
j�r��cK���Pmw��f5q�N#D>��|a��dZ�j;�8��7���o~`�UY��ue�eЊ,������B3��൵߹��m�)��(�D#��R��^RM�;�8neN�	�Ƣ�GyJ��Zk�r��093�xd��NZ͸��q�~^KqJg'^��gJ���#��=��-�8��Y!˺N� �ma�wmp2F.ӿm�d��~hT���7�UNm,�]e���ֵQʄ�j�"�1rM�-MM\~P�6Y/nx�(� ��8Lx"�%�^m7
�?��5;����d�0�뛄�+ZeH�×���sL��a|v���H�3ړFyW��[�cW^����n�YkL��xM��
2�l� ؞��!mj&d�wI�c����,z�Ӑ�R )x�۩j���RHg��"㼆�K��2���Ik\�����*[A��Bg��� �e6�2u_8�Z�Rt�pq�C�P�����]-��kj3v���ؔ>�B(�ە"��`ZT��
zp61�hC�kۨ튾 �Ub����vWU�|4 ��l�a?����ʡ��L%����Yi�"j��.����v��rTQ<cnKT�D�E�U� %�~�v{��đ;Y��´�6�<M䢷��g:.���:2���5�ﰔ���!�7��ׁ'iw��l��2��ns��u�:0���C����V�;vw��(����`���u�Xj�p�c��j��{�=�݃��r"~�D�&��}�8k��}��\�}H���i��SV�­�{��d?O��|�o�[>�v�ט���HC]��f6�|�|�?/�V��I˙Z+!���3��6<�Y4<�C �v�&��'x�Zm���%�
��,Y�l��Y����Dw&��/�����DZ5��]2{��O��ɢ-�B6�^���г��[�~Ř���-O ��ru�!�n+B��%�.��9T�,
U1&w�Vo�%ɐ>�
���wikDWsXK�!ђ��C=�jB�R�B����41h�L%���}����"I�ѝ)��n��[�x���kN��̕j7P��8����n�8X-�$���!\�eJ��!�=�3ɥ�Ec	�i��h��{1�ӷ�BLjz�Ksif��4���4�X��j�֣�&�uC��5�g�аa��~��ٓ�{C�?u�v����ڊ(&J%[�6�����
o�B��������R%\MZ}��^��:�7P�u�ڹ��(|�'� ��s�qې#Sc��=�I��ϒ�z����5�D����v:��P1�==\UԿ���eK�$�+]k�
���d]m�U��l����e)(���ٿ�ş/r!yT��L���������¶��͜.W��R�$/PަKn�H3ʃh۰��_�k ��G]�<�����Qߤ�:�A�	���](����l�Yʁ�;�(��qS�w���ǩ^��>,3nX4��r�m_ͯ�ʓ��~�be�yX�u^�Wz��)1b���s�I��U�G�`oa4[*��p�SO�S�:���C6z���Y� ��w�����mi��$�2V���_p���7�����,'�u�XM??
��E�����qQ,��ɚ2%}���!�7u���j�{��������!���*�\?�` (���"+ř��S%@3Wu6#9%�#E�z�k&�#l�I���صy��T&Mc�$��`D]H�/��<�SLY���NcA ����*�	��uJ<�����w��5�2
x�%���|i��q�ˡkQМ�4�����v�9j�&�	���Y/�8&��Ŧ�2�|����e
.��D+��ϭ�T�+|E�����CwM��bs�O{�8�ڷUn.\��M�|�iQ���cm�)�ƀ˒�c�gu<�	8�:�	�\Z�~C��#���E��5�«Uj9�"�e�+�H�6B�Z�a�v`��nFe?P�POlX
�.X�h.���� u1��ͩ����j��1����_�?�D���m�;E��D`�%&B�l�N}��	&m��R<�3�fe*5
�������UӑB�Z##�d��*�8:
w�.�7[~Ĥ�+9�;��T�M��bx��� � xL�w������wcp�_4�?*���_�|mg�E���>D��x�O�ޝ[8�a^T�x�I͖�C�C����]�F7o���7k��A��ӻw؈]�o�(�%�� �t�ov
%rM���Ac�+���{;�):���퉹�8oo�����`Ú���c���'�t�jT!����3�C�RH���{�Da%�@�4��R��S�B�Y�W���0]�U�5v!��������=�p�a�b��l��c�����̦�T�^�hn�u{�m�`�!Л	�΂`�oV;-JG�v���B�3������B3�t%���5!����W�� S��h�,�m�ZL~rAhY$],�W�F�������W��E �k}ɖ���n��h	.�ǉ���+J��g�?�U-wS݁}�^����8PY�J���ӫ�~z�+i��}�q�.��)(�5r_�Y�ʱ���}R
��.��)�o�d�8͚̉����W���؋<UI�m#��[Y{ԤDo�.mC�f�V�����C�
��H������B��_/�ؼ�Sb�xҰ��zYy�޻��!Y�<;kQNU���*a^G�嫳T�.�K��Z�=����C�4�cq��"} Ӯ\b�Lg��XVƛ!�0�>�?�NC�����2tO4� �]��W�}աl������� �� ��B��"`q/7�In�\D5�$y,:E����<s�.��1�h��;~/Q\��������??�n�|��}�����ɸ� E�I�8O3�:�l\�~�u3:a�,�����C��X�7[��6.�"�K^�;3����JkIY5��Ď��@�BOs`KvjU��|�4��Ӡ�EQ6s�k�h��e鎡�mv����e�c/]���։�l�*�w��i�'��í��}\ҥF$��I�AFLVQ\�����j�̪��:�1��?�?�7�����p�S@*!��ל�9�ӵ�-����� ����%-{HS���QTq%7�p�������E�ŗl�&_�����,j��m�.���Nq�N$9�?���݂�r���1�dکڽ~���'�.��_ �J�u��}]ɷI�:��;�:�q��#�Ќ�[*�s�5�K�O\���������n; `U犚�E��KbԸS!�ˎ�-�x�fo�[P\��͖��w@��y�3@�̅��-�m7p5�Z�~}Q���H3� Ь������n�e�X�R��f��y2�i0�N퇶��z<F�/c�\N�x��Ee�ж�c(�A�I�Q�p:-6��&�@��!�=�$��xcK�[t�_�u��B�:=�o�	�fR�IEW�6�w�'m�(0(Y9=���y̀��C߲:a��p�pw�z�	��E׷�	�2��9��r�8�٠}������~*������=L(y ,�M_?�]��*g����M�������v@��22Pl֔&�J]��;o�f4*�`,`�ګ]�A3두����v{+*ݗd`�%a}F'�vVbB�%�e�Fc�;_uƝK�h��+4O+M��R�\�
��<��-�?6*Ħ G�f�bDa�5�c�����s)��,bGȄ
i/��w����� ���W}5�(Ms9����2� AЕ-ԫa,���!?���L�N�m��U�r���M�1]5$��bV��p��i1M���d��r�;�L�ZS����3n�*K���(��B3i��˧�T�ԩMa�,���=��x}Z�Y��O��K@u���W��R*��H����Ho�H� ��^���\�E�ă&�"�س�Ȟi�PkM�q^^7>_it�[y,���`��56���d��*���+�E2X�n�6���UOyB����1��Ԧ��l�i�Sԯ����g8�v��P�x�$ل�S������KiŲ�ob���%�����;[���?��Mu.��A2�Bٱ�x�J���z�%����̲��B�P���ƌ��a[�f0�j�m�B�ە��`�,~E�s��	�����"3�q�yJ�n�~�������xѤ���@�6Ӝ�����~Y�2��4��Y��ś��*�Z�h�>M/m`�\�E_�2�.hG`3.Y�cF@-��g�d+�o?=�HQ	�ф�$�b]'����T'wK��:�؍̧��W�B���Z�owi������)Fz�����i8C,AQ֛TEA���)�\�Nhߥ.�h�� �8����.������n���_,��P?xX�4���S��`U��^>˻R�w} ��<�+/�I�iQ��ݐN��s�_�(h������h�@��;u�;�P\M���6w;��mZ�\�p.$M�:�r�T=��Z���pPKoA������B;���VHb4,Ԏn�	�g�2_u޾�(�Z"�:;�-(��N��
��:�-Og ��/|�9r���F���b��,��%�oeAbjڥ>���d��"��o�
����:���4Qr����~$�����BK��ҀIL	�31�m�&,t_Q�!+Q��F�g�aMr-S�NY����y���-gY�nث�/e�Sz�W}+t�B�ך�]��{�=\Z�+�,31z�����ɱ`U�	!O�t�Bs,F���K��0E���V�e��޽Lۻ#��b�"����;�K�>��RB�`(�մ��@���=�gD�Ώ3��!��Ջp�a���x�8�;5G��k�ˁ�6iM�J�$/�׭�U�:��	^�#I�M��M�`l4��=l����s�*I���������,s�6�b �}t�B �\�xL:ޜT���{�tL�.\��I��������I����ਦ9��'J5|hו$��CKG`Ll\��	�����c��#�nZ�.:��m%0�1I��+6��U�r�(^E���k�\�h9��f?H;1��@c"AF�Z$����"Eژ���%��ـ��m���>#-ו~*���6�;!���d0�dJy|��m5{�-�~S��6S;Q�	Wm�X�Liթ�I�j0�E��B�y%2�x��d��4o/^���*x)������r:}y������K� �6@K2ۮU[M�B���N�ʈ��9�����O��$?��V��6�Dx����[`p٪-��Ŋ������2�2 ��~�{�>�'ks�T�R���hS��gк����6�LgK���
�	�i={?�/Vg��$FԂe�m��泎��(�P1	��hp�>��e�����3@�����rsU�	��C ��ÑΖB���&���ϰ^��Y.N�'�T�c�}�X���K�m��?�|b���3Gm!ۈ�i�����8�M�L(��f����Ԥ1n],N�F����MxW��٢��],�Ža8�Y�ez��r�D�(��s���#Oj�V=�}Q��$�S06����T�Z�ȝ{�s6`�PH�Uc�x�����-�,�.݈޼
mz�Lp�n?)���t��������l��ѣ����ˮ;����E4ǜ����)�+���1�W-��"L  �i�ݴ-:#ڌvZm��c)~�,�;�-�s�p�#��qOA�W��xWa�F{*~=�?�A���!)�O���Ux�c
��l���u�w���w|5F�A�Uh�FZ�����=�e�C�x��s�9�L�5��a5IT�l�9��J&��)���\)�<j:n�)��5u��X���(U��	�pj|�s�}�3`�.BbE��;�� ]���Q$�O0{����1IC�:l�G4��'L;T���YC�̊��M��(��'�ز�<-܄�//DS�܉�����x:u��a����m�Sb�;�h����HX�~�d��=���Z�<1�}ns����#�������(��+���q�p��Wc9�C����5�*�h�]>�ꓛ�7���7�����0�A�͖��s��ʨ��I���X�t�ã�}��ͽ��i���ٛRε�n��* ��b}`�Gh�/mɈ�B�t�ǖ��F��Y�"�R���B�j�W�M	�˖��I���BKB"�w�����/���:" �|�f�Rd�%ektס��I�����I~��#ȯ�q��#ʓ����U&kH���c�.��M���@6e��1��b�=g��f��e�7��-ujyѰ��͕�̆5R�O#4��h�< �ΙJ҉�����~������������Wi&���<�?�h��������� F�v�M�:�[��&�}4���>�4��5m���(O�v"X�]�
�������mgFF^ܫr����l���ڪ"v̄�03���M���M�c���N�d(�����fő	�B;W�<�bp����֬�L���R�C��?�J�+�I�6�X��g�A�@bQ�X*|wg�*x`)�Y*�ޢ�J��|��QI���&��R�-VZ�]�.J�,B6�dT�6ت%U}Ol���dP�L}��1�9�|,E��&���67��i��[h��?峝O���?�r�ԧv�ad:i]�.�����b���2UA'�<PP��=�}�LB��j{-�H�9_�;��vj���h	�̇(�л�t���ʉ��˕�9�����l��Fk�p�_��yw�6S���u�w"���d|_�����g�����'{��Q�~������r`�
"hW����E�����ܹ�;�0dd�Ů�A��F��[��/V]I���]� ����rD���F���ݽ.A]ӗ@*��O���6�k�(�1.0Fq���_�~�F�? �L��0Q S\tQ��w& �I�ܯ�H��4�j�Q�>�*ǒiTX�����ެ��9C�DYZ�/�7h����ʲNLR�#jFʝ�����&$��$̉�+�g6f�ւ"�	�	ժ�y̤1�D��*G�K[��o,��G"+�� �(&�d�[ )��[��
&)]�o5����gE2����)v����m�4�QG�sfλ��/T��N�_%e7ɚ�t*�P���0"�&v=�I7�k�%n@��D�N�z�p��pH�͓33���qT�.�(q���'��Ξ��L�n����ެ>N�9sP��F7`>P50�����]�M\�)���U��%�}X�= �+a�O��n1�.�e��6�/ź06����dr�`�!R%+���ڱm[�Q"o��0lI
S�i��#K���N�F=X��B��x�$AfiVpz��_��k	��ʋ�u=�LVp����������u��`��L����D/��C{����/��kP$�[2>�
N��-�����^h��]��"ֵ�o_�ng��U��صǦ*p-�E�6ȭ	��%y���c,V��s4��.�G:	�p�FDsb5Vj.���8.*_�6���"������'}ٶ�"	Z��6䍻8�<�ѭ��L�L�Uo��{����k2�[��0��r�씤��1�Yd�@��Շ2A
�#��]���ť�0��ZWZ�U�o��~B�2Q��b)�����ŀ�=Jw�h�k���J�ll��q�����Ȝ]���M~�J08��[PXÃ�Amn,��I���=A�µ�ؠ�O՞�1�����^��`֗�;��@h�!���I�d1����#;&gn�)\���y��SP�E>�X+W���Y��f��#��;/j�[��J��� w�!�L�q�����,�Ȳ����M�F f�-�8\3m���j	��Q�!�쟧|���Is�SO)Bď����5M��Zl����2��8�ґ�E<Cд�!���`M2,uM��9'��h�\���K�)�+Յ��@
K#qג����ј#���#-q�u�4Ǘ�{?n;z���M&�+?kj���B+޻�I��[?l�=��6���7�j���
Tڟ���pq�,[@���
�v	�������$�NﳼEٍ�)z܅~�		�Jb��^�v�}-6�`�#�>��o�ԁ���^�ǢH�Wf*�RgN�}�9)�]z�������_Џ2um��֮o������� DlW<#�����+�	(�RNR(�Ӷ�7��7�vo�]���˷�;wc��ϧ#E~aR�{7��B�>�,�ӌ��*5lQW:BSh���ac������2/ �Ր�Qr[��2#�!y��*Cq�"���O�4V��N�ѐ�C+�O�C]<��[Y� O��#�v�ъ����g�+�� �Ȭrl>O&�4_T�7P�^��ie��@�E =5�)��'�D4�,D�f_n�J������r�Ǡ��$��ĴSY������݌�
���bo�	i���J8��i�Vz~�L.�f���P.� �,ǁ"m������:��Ȟ�@m@��&dDTz�sh)0�8�kr�uk��ˊ��TF7�EK������R�׋����=ݻ�?�2����zH'��u������T�A���Ԁ�Ʈ����~=����p�9r��O䐵���؋M��(��]�B���8~�D
p��Kh>Ή%����a�r�ת	ͅ �n�����}x6f�M��GI���c�޽)F��T��[Χ�T�`e���zj]�	'.�j����q�y�g4=%�`qD���_�ӵ؋G�l�@71�$���Ƴ�m
�|2���h�$���p�X����}ɍ�]�b������3�z'��=�Lîw�F�֒,.�vEE�Ìz�g��jj�,��G�tn��D��g*=�8F�P�}Zs=�"7��E|�p��[�;4��i�m�3ѝ�p����� >���@��v����zZ�c^*oc��K��96���+�D�?vS=���b0Dx_���
�{jxpJ���g�غ���0Q7��E�+���-���p&�YО�%�%v!#8b��r4t:80���q�pOP��8y������"e��]+ rvt0����e�K>Yd&����,�G���y�~>�v�a�%ӊ<���� �������sٻ��1�9��fGQ;����cz�P�w�U�}��1��u��E����T�˦Q��1mH���y���Ъ�0��m*ɂ�b�)s�c��H�i�`6|��0���S� ����)�^�=�a��$Y��ŵ��6h�Чg�?*g���u�pA��ڤP�q����7sa�iE  ���a��P��X2,j�QIT�-��V@��<xE���R��ڞ�u),o���S��H�G�^�H�=q�wP�� m3T�nV�ΐ��#!=~5�۴���&|��τ ��pW�E�C�����JWt �i��z��1��2� ��̐�6&�(>��mh����S��]m$EWڏӶDh�X�|��P#z��I����9����_U��-�L�.����Ur��=��1Z��=3�rz���Z�ꮣ����P�\J�
�b�[�IO�ީ�i��R�С���ɛ]vۇ��)�2 6_0�<A�QΞ���T�`G�m3�9�(��G�tW��d6+۰q�[�U���+��Ʋ_t�� F����<��L�ɤ�u7����sB����*�gs�Pb�$"�́,�Y���Q�N|,�\0���2��Z?L�%"��/��N��0(��fM�6�-|�`5�u��3�p���|VVDϋ���W}�V����BO�U}�� �W"��&���+�nw}l���*��{y����'�ޮ�z��q^5���ͷ�|y�)O�ȃ���[�֛��l#C/���Y���6�&m��5��x2�>��iRV"^��h9sj}��Ŗ��f���
lfy�W�r�pv]Y��1������}̛����~��2?uR6͸;6_�涝 {�/�Κ��VH6�^��%.�Q���Z3�8�7Ĭ��$`��IK��u�W���U��r*n��;���E�*I������ϥ9z����gU���o�оR2x	�1���C�����R��_�Ia��V(G���ޠ�V�6I����u������i"�:�#�Y��TZ5k�dyqv_Qꥎu��)���,@�;c����,#po���I{���x��`=m�yv��8^jlE@:O�r$N�`{�l�wϮ1O�6l�oWXc��vhX �����
�ճ��FN�߁dIJ' �Ս�����&�0ʃ:&2�}����t�u�%zf��ʉ��W����υ���Wy�@��1�~��5�5-6������
���4�",8�&
�J��n�:�\9Iط�"K���3��A���PHuے����z��a�m���=7�ۺ��z�[��X^�q�~S�bw�6Ҭ��גx�R���=|�h�}+@ Tc*y���9��	ӓU�$���>UD^
Kd��%c��?a�-'g����L6��j�@��Q�� ��d������L�����A%t�-�q����9߯� Ư,1.��Jo�Q	V���1��ŖI:XF�T�>VA���P;5T�@�$:���ZoB �0�@�0*Q��D�lQ���.�E� 4��Jf:�+x	?)u)� e�M�#p���0)E�?;$�+x䃳*�p�+�/�j��b�Ma�)�q�ʁL�-��ɁZ�#�h�B=��2z�0����5�º�&G��w^����>.Q���+ᄀb�U�L��F��+���U��m�����+ĺ]~�Ϙ�dk�{ٻ��͘?�՟�@G�T�#�s�~��͒�yNhԧ�%���(��:'��>5>QN��B�q^��F=";�Vn� @?`�iu�	�(���?�����pD:�:��P�jہ[����>��*9AMc�ª�&�TϾW8�*��s��q$^ŪUr�.�_��e����ϲ6���_}ú�G)A�Ek�ɓ��BY�0�*u_Q,�s"�# ��!r���`$}4^Nɖ�'^�q��r�_�,�d%�V-�Q�\�]��f�' q"7�V��^/���hÎ��Bڨ���CDy�Y:ο�H��A��ً0��E�V��P�����N8  v�k�I�&��"��w=�[1�횃6�^�eｴ�ں#�t2*�j�B'jŋd
Ⱦ�uB���Z���A>Q7(�.��A��1^P��eU�BNId��I<a�i����m'�|�Y�9�PW���nd�����j.���P6�!4��^�%:*{�:w,{�)^��I��V��#5I�wU�� �A)�=� ��~<	�(#d�f��[��Ky�5`�봊�㱳�Ϗ�xf�K���s+����Q�?gk��h�u-9�����z���E��˟����I��x���^�1�E�<���qJ��1�1�]h�Ɯ3S38��3�^��V������5X��u�	�4��aFr������3��P��Ɇ�ҧ��}�e�� �H�F�9��]����Nd<���^������M>E��՗h��>Ή.X֙T0�k�V�с���sL��s�cOť�w"�Y�CjQ�V��m� u�Iyd5�/�4M\���u��+K���-�^%�9�a�����ʿ8�2a�䢇�-ygW�/��V\b9����.���w@
��� �J6�HЄqFn�!Ѵ�ySW��sx�}l�O��-?� ��p�d��DL"���x��V�����Ӆ2��#����:SYdx롢�ʆu?��ztlsâQ)����yQ�1t�;j��\��1>HoTi"6pQЈ�?	����=1E�]��y�"��M�����\���E�óK����C3�U2D���D��C/�ֱ�0e��pM+��-w��2�u�q�x���u&gg��c�SX��*6�<�/���m�5�A|X�-�'�k�(��� ��G)�Ŏ)��+�)H1��$�%�R+!�L�afP�+�c�������i��!��6�v�Mtyh
��Y)��F��y�P2�=�zY�w;��y�`Y�F��}��D���u�x�����:	mTۣ�C��2��M(�Z2p+����k�%���KX���6�a�(d��F1X9�ERH;��O��V�����S'�Gҏؙ��2 ��T������(̰��jd��]�E�⟴�YG��@��G�"�2�[u=^;� ���a��o�8�'��O�.G$��48�V�L
| /�"xvW�,C<Ca�O}h�Ɓ+.�n�/kX�*E�?f8���1Q:���jϬ��F�5�l��ͽgߕ�T�˛�YS$�]3I���0�Q1	�bL`�W� 1̤U���Z�蓼��)��	u�Ss
���e�E>��ݒ��5Z����lw([J����"�j�=�f����N�KFt#��P5k
�ƅ�ї����-'��/6�T�&}���%���9�jݱ�+��O�b=��?����"B��['	�pS����O?R���|� *��B��;��_G$g$��< �	���-�ОxW[~6��_�:��t�~�@a��yfS��b�~�v
&_��j|���+zz
y+]P2�	��l�2ڱ}�f~Rd�n��F�/���%��>�;�BsNg��xZ��k��˰M���G�u���N-8�?
e�LM���&�"ҏ �=%m���(�n�<�Tߏ�g.\j]�Xk�Y�f"f0�����dbi�G?�4�,��-Q�2�w�?������E6���T�y=Fn|�b-��sBН-���xW���b�_�N�:K�vy�!m3��CW��#��N�
�\	
�%� ~sYWp*�m�r�n�$�r�W:x��&(J�������?����̂����(���[�j��k���z�u���/}�J^�1rq����Y\C˚��G��-$�. �7��﬈��L�T��I$�T������!��Ph�'��`e\e���a���lWzj�ݿ�İV�6X_ �d�W[��oT>J��;�a�!�0,��QP?w���U�%����8��I�0�,熗��S�< ��?lQT����[��k{��.��&�[��d�5�Wp�+=x't.}8*��J,d� ��r���-o��V����s�(`��d�2JVr�^H�����������o�R��܀�݄���Z�)��6�
��ϲ"��*#h�-��� q��+a���sٟ����3���.���"n�Ο���i����]Wl��^>�٣2ً E��=�~�f��)'7���)��qo�wL��Hz=@4��..b��lC����>R��ݕ���B;�s��*���+Jl�ɖ��db9{����d�'ۓ���$]	&>q4cCS��R�[.V�r�Ox�}���t?\��I_&�����y�ʉ��O�l�%���Fh>ent�y6a�Z��D������~N��7:?�%N,��4�N>�!�2�c��80w;��stV��͋����_�.�Zƽ���Q$Q{�LV�<�V�"�h��w�I����f_Z�8i�eԎn��:f���+qk���ϲ�ŹPyE.)��d��]6v���*��ԓ�/��q�VA�nP��ܛ�Ȅ���Xe��)�cR����+��-��"G'5���r\j�ub|���z�/T�T�����n
�~4Z{�
�3�$O@2�Z�֦��:���,�D#�����%x�z{��<�?œ��Iϯ�V����� Z������B�	uU�@m�hc��W��
�(f^=�\����*W���hC��C��TrVxʱI�m���D�a�挹���ڧ`;�|�1\12����E��Ƕ�Z�b��OB����Z`��ff�Zss!��7
�3���M�;�wo �gƵFءC�$�n^������<�ʜ�v832)k��>̄�'�Z�������%���3 �Ւ �-� �0n܎��`�v�N��遬�݉���'�֋��_�cԅ*tP��ã��s"`bv4�\z�;��i�
Y�'o�TK����b\��u�te�Zq�$ĖB ��Y��rژ�_����C�T-�Wy)L��b;֖��6��a沁�t�h�� �}��?|�&� ��$^~��-9�h+��y
S��O������kٯ���Q�
@I��6�6x&X�����{a��z�/�ymGr���a�s��R��I(0&�~��+���)�+Z�⥘�Q���>��H,�����%m�p��Ɩq�V�o�^��L�䠥k�$�3:�$3��t���� E�o���F3|�&�G��$��+4�w� 	����-h^�W�}����:UL�n�d"@)���o���w;�j�� <�`�3i;��I+�o
*[�ݲ�VSE��SRN��D���O�R:'�Ϣ�a*Ѡ�a<iW��q��$��J��Zb�#�g��l�ƔF�����)���+S�4�J0m��w�Ӓĕ�
�b�=�rv�+���Τ�������O���*��M�9h�u��g����垒}?�PJ�1˙����_�a����K�.\��홍^L��v�x ���л���}��
E]���m7��K�b�_D��(Aǃ3gD�/�c(�C��rs U���(��t>���Th+�j�!$G$�Y�!ڙ �-[S0;��l��;�JI��ζ['��c&�vmF�@#��̤]��}�`�� �g�`��*��E&P��A�͘e�!��c���*�_r�i�@B�D��$�1�2C_�"~�>I*�ٿ"z�ϊI6_�?�O���+�� f���yX=��Җޞ6���
 �����"g���K�R�o���K���i軒}���}��>��M0���
�B��m�DAJ���6��Iᅓ�p������v��MR���U��h�Q�o� �q�c' ��r��������)�����Q&��e�b�����.�,�H�mP2U�E"w���6���m�$���g7Y���f_w|�C5�Gi+0�O�b9�Jv_bK�����忶�U5�L6i���r@z�K��ڏO�\�W'ڐNT?��&p�#{'�ǋ���d*�X�SS%?����Jm^E=]3[��w|�I e7��}��'�o�!����9MxT��B�5�s� ��mlk�>d�nJv�����w�@�U�������f?+Y����C�sMF9�8w����sHCN��5!RL�q�Ѧ�\S�g�v�_�s���ʽ#e/.l���HC��H��`��9�.r�+��P�v[�#]��^N<̳�*Q���m^p�~��:1�K�����D�a���3����}��5.�}���{�\,�9���W;�U��S���l����3�'���~�N���'~/vq;��}Y�竹^D"Š<�&�&�h���i��b�$������	s��b@�r�mJ��TV����ɍБ2|��"���(ms���l�s������'��b="��?�I_��QA��id�2H(?�s��������q�ȓ�� ح��-M*�K�I!�y���2�[�l���Ѽ�`��AgH���@�j��?3����3�!'}����*b����M�� ���BW��4g4#0�ǘ}7���
v���/8!0�s]
�4�71��0&gm���U���{i����S����D��q��KS��zw�ҩ!>^O�GΆ�k���`���p�D7afP������Ҡ}g2Y���$e<?Pz���Wo{���m��~嶈@ʶw��c�+|OH�Ŋ�j� S@,~'f���#���F�jD��m�V�U��%�5R�b��,?�Q~~�G9��#���{��|2�-@$�4>{� :l�+����l��˟�ć�6�V�eǍ���+Km�C����H�F�xS�ug0�^�I3/�����@�q4Vߡ��ښ���c�nX�4+��M,�Ӑcc�ddn���<Y�=&[C�B�J�`�6mM������G'�)��L���������R����euS+�m]/�.,D�P�d��ڢ���D=��!��Ai���T����,xMU�$��'m#�tkV��)�8��?�H$<��5���;)��V��D�@�B5��v����|z�"�`6�nov	 i�
�7���X���a�C�h]�� -�H7�TQ�~�Ĵ�i�}��N-R����
Տ����F~�7-�-���p?u�����fIi}�^�Y �{��0�F�u�t�"4��p���p���z�*�9�ﾋ��j���	�cw\ȏ\�P��EףO��� a�H�V��D��PM��utiO�܅���Լy9=3���W���:*`�nOK;�W�!��@�|Ѡ�b;=����ΰ�\�R5LO��5wf�<lT�w0J���ΑC
��5��X�T�E
�-N@:�R���q��"�T��vr����Ժa�炩�uW��[0谺��!J�yX�:��ڀ^E11Պ�KHSw��E�j9o��"��G	��/�"f���'�yr�� ��k@��P�X��z���LvF�F�%e��I�s���Ne8�>2=�t�JJp(�j�L�ՊL6�H����%�a^��<���qN��L��	�u<���Bd.�'�jm��|�|���P�P���H���tH�$�)��	 �h�!��J�Ũ���Б��K�i�������W�]Ff��J�j��~1��lF?�����3dτ�?����ԑ�s%s�g^2jV(�#ʾ�V�z���=��S�����	n-���S���ױ��S ��B/����\4X�$5]�"�{́ڍQ�$�ox������7Ht��}�N�.��t�#���Q)�a�(mKws4�,���`�F�8�'��d0_
���-,ֿ������Rd�7"���.�B��-X�2m��%�"g��Ҷ�����*����Z��[����Rsـ���tsܶh_-��8[/�Zo�t�$�r�p@3��6o�Uڍ��mL�$�{��4��+h<�5.Śm���@����4�CfL�=�c�����)ӡ�cl����M���s�	Nx�9T�;{`��yKُr@}�[��盙m�tCSm�Q���r^ds�W�+���Zw7T�o<�O2���{�k u�E��&G�W@�g���KUvs��>j��K9�=%�R�_ʩ9�`(@�b�6��нڼLF���M}(Y]YV|� �awx*�Y,�]TX����p�y�n���]�u�Ln=[ᣳ�y~��7D0఍f�	��y�U�I�^!�߾7�սз�	o;S��#p�G�rF���n�{I<吱��ҽCi�)7ŧ��I:�|F�X�?g-�k`rL��a֫	t'y=K�c z�9��~@�s-����+��?���H�\��~g��8�U�LU&	8Wq�J��J\<k9�������ﱜ�9�nw3���h ��/H����.�J�7����si��p����3�N��X���˪y�HL�I�m�iZ۟Zru�$;"�g�V�S1M�gR��OS�+��\]��R�n����k�i�x��ck�v���DOZ�OG�̕�i�����(@��Ժ�.zX8��n��l��Q�a<�E��&z��?��?�}�	F��6��o���`{�@v���2�/ڬA�Z�@�\(����8�P���,Ra���W��4�G�A*@-���D7����[
٧X��#n�!��k>��H/�X3M1f�h�Ca�Q���3���YgL{�5\r`�f���*���QB�^���9�87�)ǌ+�U�*��f�c�.�+���i���_�,ڄ؇BQ�u�#��d�W�暠�K��{�%��x@�R�}��r�\��%y�U�=p��,�HZH�<��w��'K
�$,Eכ�D}�Ł��n��]�'�w����5�׸��d� ���l��	��ݰ��z߈�H��#I�l{�B��噺s�1�vx��z��$�o��>� 5H^��})�o���;w����IUO��EQɍ�l��aϩ���;�^F&�?��U-,�=jm�곬�z���)�^��n�)X�����Y��0�۝�����-#���c�~A,Ȟ4X#�䘗�G��l��{��l�tS��'?fs&�9��)gx�#��шŦ,���,���H��`�Gl;��F�t�Ƣ5�? u�ǯ����B�\�����b�z �u^-��P�p�eD��g�Y5��C���5'�+]6�?�OiiqC�Z Y ߪ�`ס@�T�7qV�=,��!�B9i�����Nf��9IU��s���"�4��(��47��qG�>�������p����=U��p���޸5�x��kI �� 1jd�g��޼*���c�Õ�3�y�n��U"U�>�z�of���%��I�l�6l~$B&P!Z��R�6v��:��H$W��Mw�������-�!_���l�������ۣ�d����N��W��B@d�$b���w;Wd��E�4�;��XD1כ���e>���X���	\�o(��V:�q?DV{�#Փ���|�u,��;�~�ۻ���t]R�� rp�����̍5+���S�_�Tԛ��ԓ"&M�T�j�]��?�.%�|�\e`:�oT�N�)���}-��x��D�j�����Q�iف-g&���U��lV ~�r$%�=2 ���cKn>���� �R� %͛�[2����Ҟ�~ ���ZY�Ҫf�	��SsQ*V���zN
���1�h��A	�1g`uu�
��tę,"S��`�>�[���J:E�M�S��P�/���oZ|ܞ�O}�U�O���^u��a�74	Î��{�~u���ORvl��a��lL)�l���~�bGo�,����٤�0�:�y��I�~��8��	�f���谲bX�ٶ�����G9�g��M@-���)򇴀�,�>G���������Ȥv�'�!oM2H_L�N�.N_^�#&G�?RF��ڸ����h������3C��&.���J3�f��R��f|�q���7JѱW��]���^H��b�lD�9X%��$6��%�8@}״��5�˰��D4�������&Yړ���Z<�wY�T�kj6���$\쌿k��7��e.�5�V���"��̭�7h�<�Y���)��ܜ��%G�1�zNm��A=å���r���CR�!���W�����[�H���c49\&�z�x�v�'0RF~�/wP4ڷ)u�o�lwtv�",�C յ�ʾy�;3�������)�� �����B�ȋ����yW��LC��~���n>��mɱz�b�7;�!���\^J8?Ch��� �7�ťf�g��9k�=�����Og��ay�fG�5���'�xL������(�*S� ʍ�|��H�n���ytO�Y�E��Zk�����&ᄤ���gK��]�2��
��K^�S��CДсJ�g����Ա!�)��ǵh��HD���:�6�i<�^a8�(��Բ0p�i3^h�/tq�Y$υ/��x@f��ޘH�/�f�(��a`C�� �Ӏ�c��z�^Fs)�R.i_����������d�tg��ز�3���5z�Ʒ}�P�m�!Y8���O2��jH-��MIV����bU��cs��Kۢ=��$B�8�U�ř��bW��p(tC>/C����9��͠�D7w.�U��Hp������Z9�	'�5�`����ޜD�'h��/�K�����Ϩ>*gk���"a��:�}���$Z��@�&��R�&8�����\�tfE���*�����?�l�-TD4�9�R|*ᩋ�H��o�˥���
�}@h�Xk�w;�&�����
��6�Q���`0�vO�� [��d,OV��%Ҧx�Z'ګ���f��V�\TIdδP���'5��j���^ʦN�#8(�Ti+R�F�o�R�;
�$0!�X5E�%`7�-C�l�M� ��#q&�.|̫Yd�������'�VL�cN���Z=^ֻo��JƤ��䤫?��T���꠯����j�$$K���D�Rl�fv��Ñ�@�%�%�q��`4!��H�36�G ��.�@zV���A���e,B���P���YΙ@�Ѥ�r���l�eV����9:6���ɏ����=���Pgl�;��ژ��A�;- ~)��	����N��O��$�ve��2S����+�N���Է������XECu�.�8����-�� ;���zs�<:�`��E-�ذ)@x�ӆA^��דL~���Ƃ�����ͻ�?�ӝ�������4.�Mh�Tp�ϱ����x���f.�̆f6�_42��]���>r��C�J�T񞡖��8�A�l��O�o7�f�qF�-�gAK��i�I�����ybԻ�����ҿ�ĩ�Ƃ�m�O5��6Q�H�����O�W�ʈ�\C�4�^��/d�ё�� 7��؄F�H��?��JZ\�G�s��)6��.��h���jy���g�v#���}�(~��Z�]�)|���ŉ��D�K�>�-����}�\ 1r�G#�gDֲZ��ȏ��4�:*�94f���^�ī�\�� ��P��^�%{Z�EU>5��q�c�*_d��oqF���x��A8�jRO�J���®V�%d��"gc��K�a]����t�lv33���+0p|�@	\��Kv�m�3�\U��.��K�+�����(�3���.����S���*��6�T闒#4} �RԀ�E;"��ffg�G�>n]�A@�v�$�R�Y�0��Ah���ХN$��>&s�������D"�ig6R��>,e|d�nbӤC5Nk��L!/'�@� \g�}�6�������*K ���k�F9*$پ����G0a�_��w&/�1�h?�J�8Dp�iT�uz_�K��� ʺaG�����G9��+��KW'�8э+�����Aw�~��!�a�;,N�K���>���O9�&pMY�����/+Txk��J��Lߖ�:�@��'��'���A�kH&3ݙ���t�)�޹�"'��|�L�=�U���T-}7�YK���W���P�ߠ�t�����Nr,�P�'=��%��3w
<�����L��� p��W:xh�SUt;�9���a&�P�
�J5��VF~J�%��<[t a�T�%D�R��?��}����*l����8�/�2@J��<ã�+�>/��@_��ەD`�>$��_#�PcG/�WK���;�l�C�;4/Y/P��'��]��Y�7�3��[�#+���9��Ɇ�2g"0'!��ϣl��{!�s��?V�óEJg���y�y�z�$����w�NJD+eg��3�A G�����I�������'���M�
W�2��#��'e��9�j�Of'�H����ۮ����7��Ԡ��:���NO6h��5i��P�J~%����~ŭ�4]b��"��85/�������_-�o�m��������7����@�_k����01�b�� ����;lm��;�������e�o�)~<Ejq���{F�Oٙ�X� ���s���?ʟn��X�� ��DbH����F�;^)�^u]*c��-{?v�a�-��}-�>��k�'�L��N"Y%N	*��`�g�p��A�4���l�=�TS�#�"��0�xE�l�N�ct㾍�k	H/F�am#�9�'��ZOw;��Zd���#V��y�Z(+k��/9���;�Sz߿s�N��q�۸�9�)t���M�c���-���a�S5���5����TC��9���M���?�@s�2������A��d�\ɡ7u��
wo�z�<�9Y����D:
�{5U4j�pQ�jP���d�Ϊ��e��.ҧaCJz9*&-���+$Q�հ��p���#ڹ)v�6*(+���|a���>lU�YUV.q��V����p�惼� #��ߋ�{��9Z�54�+\���i"%�\�&ٕ�R�*�Z�[�6��G����e=��!�`�(/X��o��J����f���p�=�F/r^K=��R�O��ʣ�Y��J�!��Q+׿��ⳋ ���\��}Q��N%�Q��������%4U�c�����M�3/�~l��e�m�`Uz��������F�Mƪ�����3�[� k���̣�s��tI+0�ϣ��1 ���&�Q_���/�#\婍��Dus��W���H�+'ΐ�|g1n1uo��p3t5d��&��l�8��� �+;�`��y:����c�����q�/�ts*]��ks�l�a�^R���H*{�xLqʵ�b�Wb,[E����Dy�5Q�u�@�	+}	�)j�q�cB�;�������24O	h�ݾ)y��ז����:| ��~S0�3�8���J��πz�O�� �K�W�؇H��/(dΖ���DcB�MAH�$�p}����J!�=^&B���;��H���D�d��ͧ��l03�=����O[Wq�ۼ�,����I�AF�����X諀�d2Ɔ�5�i���߷׆ks��2�Щm��~`w�֓�l�;�W�n5���U�$'^�֌���[��2��dņVu��qtX��P��7z�I�G�q@Uω�w�C���v!�ۏ�R�I�'�N5^��4ZN6���xQ+�g	�}i�TUQ��/ �~C޲�l[ٙ�F>�jKj6�V�ځ�$�Z��B$���
�4�H��5;0��̐f����*�N���ǝ��A"]\�ۅ@/mL��C�'�P>���_=�\�za"j�$
 �_��J1��]�&9���@IT�}�^��+��om!u���$�_���-$�~��#�%.�
4�}e�7:,�ƾ�J(����+n��� \�S��B�����|R p�qv~�Bȡ�z��.o�����`�0��������ͅ�½M��%"/�]+z+K�S�5�;�ddj*����O0�9I��e�fȸ<|���(ﾄ,)�����K�ݦ���x�5�ς��)���\�t&X}܀:1.�DL�;���1'�����x��pH]W���w#|g@���dt^觳��U�F��6�gyn���8hAg?�P�8"�A� Iz|���k�7��Uf։���y�f�[--�y�P+P�D=W�>�0i�Y�m.a��g��套��^@�?�󓭳��I�����x���[Ğ�Z���ؽ���G�76BX7tE��I��T�hH��B��)H��Q��(�4�w�p:�
��g*��g��lR�3BҢ�ppT�c���r�y�+���f�bY��c4K�#8�> j�:�d��&�<�3����n�������Oz@�`���Wp7t�^�kV{���7������YA����=߁i�m�r���{;$�a0�<��XF��e���0�ϖ�7y!�0Y�2�8�u���)�W��lg���g����|�A
D����{-�9\ZE}R2��4*�	�@Jnd��k�7)k
�w��v�`�
s=����OZ�R4�%`�bg��^O=�N�3+~��w�c��<�N�z�%�Z�=�����rۋ͇�`_������;����(�1� �������]ǒ�l��^V-j0�UO�RW���Ӹ�	��r���%�E�;"�7�bީ&�6͖aL� &���)�-ג�rH�>Z��#������!ZgrM�����!걫MqW aNqK��ho8����C'��L���%`W����S)BI�c�U�m��E\�C�.:9���I7�
is�t���0t_HҺ~��3��tm8'�����!]�W~�yP�@8D4�lQ�=�� ��^*>݇@�E0�(� |�蒞���\�I��b�BL�슑�&yj� �H��K��V���BC�e�d�B٘�NN��\2Y�g'Vh������I��$�8ruڠ��ʣ��-�o��x������Df�:|Ǫ�ׯ�1�x"\G��>�B�M?_Qt���%K���#A����:vnj��'�v7E��b^�j<7[�� ��D��\� ��F��qȂv�tH��s����Q#.�v�Q�����(��v��b�P�q��U�,;�FL���K@�'z�i��H�,��c���pY�M:�+g�?��	�T�y)�2���n\��5s�i9f�~dHl��U͙�G��	��h��=�2��pY��´�߶�C�P��K��m�Umxh��%�|P��;wx2�[����<���w���,�Q.���E�'+��E�_�	b�H�Vw�(�@��Le�`dB���)�^D��!�������9�z�j��@���v��dr��D\�l.������7|���Z��}���3�j����SD�җ~�1����F��.$���E/-J꼉����2)�`�J pa�E�e�̲$	ʜ�U?(u#/�S��c0��.���e�UK����;k t�K��&�A��GQ�c�SH���g����s�b(����|��gI�:�!%�֪���o	Z�?�)��_�j��o��iŜ������&����mqE4q/���Hq�r�g	*-��&B^��t�]�efvҗbTG9r���"9�{�(��QE`B*��eW�º?R�� p��6�?�B�r�Y�p,�x�˳��t��U�-v�@?3����F~T��V�X!��w�i��]�V�OZ�)$��EO�SA}�\_���?�C���Uw����2M��$F%�hjR?���cM���������]}Ȏ��S�[�p���,�H�,�Dm	�o�:��[;���mџ�8�q�Ϋ��f�e
j��Z"�rV'��_wc�PC,�BLF�A)q�#��&����E��<�<�o��)�2��p�%��z�����S�szR��S�"tZ*�"]�̓�&� ���O��i��
�XX}L;�Уd�9��d�K,����Lӈ��'�1�=J N�5U15+]Ǉ
X!L�a=Z��%���� �嫱[E�<���<�b�Џ	����Ll���Kk�IÝ	3o\ �>=1������e/ۺ�7Lþ�J=�S�wC&�&��"�\��To�5x�����k���;�T�9~�x@ӕ�?gs�������F��n�\��.Ct��[s n�r��J65͞}'��h�$�?{�>
�2�R��|7$Y7QNN��ry�I<�D]��E�ǂ����c���^�����m�i������"ig�r��틺��ӛ_��p�$�~��q�u�0P��5��|��*����q����� �B �:� ��*g>K�P��r�����p��1���9ꌒq��s��� � ��/ꤺ<��w2����4sHH�ǻ W'I����-5%v5�]I��	�j��'��o`��H�����HO��8˙㪢�޿5d[�E�`�5>�}�M��p\q�T��1�ه�� ���������:}Bi�2^�y��g�[q��LL��b�����A=F=49n���cq�`+����݊�G)����1,झ����7���ZR"�F��=�m�휧����4xr��Q�a1&��i|�aת�ȉ�.��JJOd�fe�(������Y8�� �?�-㎝�B����l��zSaD��+M��p����!�|y��b�Kݡ�^�$s���3WY��0H��� ދ�'!k�[1{�$p,7�]��5R���6��X�]Ưa¶�6�Xx��B،�̦���Jp�������,���� �Yy(#�2������"����B��b�������X��$#��d�aLc����#���J<u�-K�5�L��(�)���j�	˸��ҡ��i��.L�߀g��Gُf�W]�J���H$c2�z�;���֪��#|�u�$��¸64���������<�E�M��y���M*��^B���0��LkvW'�����>	��@R�I��wq��5���)��)q窖�fU�בc�Q���kk���LI��Ņ ��N�J9&��(vtQ��VQ]��X�LU�[d�XR���W%�ʜɌ��O�ʂc *�o���W��|� w�t�%��p�b����#k�� �}
}0����15^b<aم&D%JW
�9��h��\[�5hUn�Ğ���q����� Ne��{�v�|��V�F���Kј$�	f"�znP��yBP���*�4��N�j��,��>�A
�������y\�}�^��<�{��#�c��j�E�YV.7�ʌ�j���x�+ש��؈_�� ��5�����{�h�#�{1�;N�>@R6�5λ�)Mf������!c=�Z��!;��u�S�L^��ZK� V��q��d�f�N�߇#���	3����h��Ŵ+RrA��;�J]lxaK�a�I}ۑ^�,�i�p�UzEW���TJ�v�\��ă�0���Pу��H�q�4o��ёOfв�������t^p�tk�vsrۭ�����۽>e��>�x���I��H~����)x�g��
�%FmxQ�#N����Pa���J��9�G�(O ���4��L-� P�~�BM0���ϕ���������\��`af�$��Kg��(��ST�+՜���Baz�y���h�<d�Z�]�^D����X�վ���S���uI�]J�.9�M_zƢ��ޫ<�=�g.p�8� B��t�6<~������YB�q��祈�i�T��Yï@ ��1��N�j�=}&���E���] ���H��"��cT�-zy�#I���}�f���3�Q�1�-7�����z_̢�� ��]��G0����}2�j㾝_*�Mr.#'�B��0�Vr�? �,��Tʸ�
\�缹{ h	�bq��J2�<	uTy��v�\��gT!w {Č���6������+��^�-�ޟM�<G���x�Ҽİ4� T�i[�yZ�`�r��d釕t-�2V2��d�!Xv��L.�F�x|9&0Ep$�IT�ߠ��L��`ڹ��)lI�Be��gbZ��g^��Z�Y�Lh��Ͳ�K	�\��m�2<�
�疉�b�����m���u+�ĕ۳a����=���,�}�k#����n�;�����`HV�b�7���8H�;9m�d�^�הAEEbe,���Q��[�/|�{1fh�9�u���O\a/c�[�#����\q��H(����/{��]u� �F$��Ѷ���V����;�;�G �H��B��\������+3��g���n��,{�"������)Q��Z���e�"\ȯ�ot�t4i	�������"�[v#�%o\����p��u۹���F9Ԙީ˧%�Xe��D3Mʪ�/y�l�ᦆz���&�v'�<����Z�^���pf7����R�1_��j�3��MTkI�}�]<�׎�Jw��s�[H�R�%�́)���q���V�����z:
O?������@�R5,�+7~]�|�}���E�b��R�b:��m��.v
���Cm-г���L0<d#3tC:>Sn���ًa��v��'��qٚ�m;�'4���p��)�r�l��A�}R�]S����?�ܛc�������6k���W�U5M�� UTCH���E��%F��c�j����5&�W�"� )Іπѯ��N�[:�̖h�2<��H�-�2��'�;5�$�hq��L�>Ebp�Y%�� �t�ڦ�EUR�a-�S�FG��3�/�mz�1?
�B+�gz9�v��ͤ�2�򭉋hR�֯�J�H ���軭^7�w^�nu�"���l����&��隂��㸹�YH����F�Ct(�w�݁"�#{���͂W�fD��r]A�/����e�*�(@C��4��H!C�5�|ׯGƼ�z�$���%I��B���h�QC�0���]��g������+M���N����+z��P+�z��韁��r�x� n��#]�ӥ���p�T v��qG3~K����R�	���1�$�JRP�b�]#�h�W>�a�kȢ�;O{�Ga��L�V"}���{�1�S[����H-N�B|��(cA���J4Uk��F!魳�vO%�3���V�Nڪ7�'%�իkd�y�{�����)�������c;�<�o�o�-��3�� �hܞ���d:c�}r;�kz�5m�*4��gg &�Xō���˶�cߤ���RuЛ�^��	ӥ.O��4����<i���|5��饄�UA.��->���E�x'h��)�q@�ރ���2��6�2�(�#|�-/W��/OG��?��r��G#F��<�|z����k�qӑfxU��ΰ�������9��z8�w2�֘:�� ?͢"�-�F�,s��J��wA$%"o��W��)�����+J�%�v	��E���wX;���'<��/�A/��\�����f�Ҷc�T�g8�&�����*&:r�d��;�G�7���.W��S{�tP��8^苏�;'?Z�*���}���:�K�י1��&���V���tʘ͚�b:w�[E���?j������)�ݽy�;S���>�@1w�<�����������Aq�"� �c��y�3k�aV2�p��'q���^hd�Uj�L���S���c|�`���pF1�����1ls�l����M���>a�LN�3!���X��뮽uiu�x:ӥz �ɇ�vO����\~q⽜^5�F�U��1�A%�+z�@.ȡ��u�=�/<����fg��9v�ӳu�z�u���;z�v�G��ϺG�h[t���T흜V{gl�g�7��q�=��3c �w�]~�a3�x��,~����Gi|m�wY;�+�޾O�#��:���jp$-�_ci=���Nbi�U�Y�&�����֚+;��"q��&.1{�+V+b����ե�e.բ�1��(<�S��+a\�� te�(�}5h&�Hf�(�p6��s
׹��e'�Xd��\��}Hn��t&�E킐��'M�����p��ΕC`S�Ru�֗<.��ߍx��=V�nTXƴU:��ӆ��5W�\��Zlp�lTULk3�Дu\�0L!�nX6�?K���EA���D:lX����+�`6�K����J\�J�r��r��=������N����>�5�"ks���8N��[��ԤFV�>�.@��/��}�Ĩ��ϛ���g3eL� 7���X�Iz�>���aj��G*�R= �633P�~;��>?��I�W�-�����Bu�߮Y�=��Dzyi\��K'�7e����y�L�
�&)SI�UM�E��V(F�48,���;�4���AJ19��^��qC�������$��Ĺ�2ۨU󦾱���/H�{�k��\�e��Vs8�]��x��Xf}Y�d˹�և���LЛ�f�[Z8w���~ϒ�X���-F���c���1{�؊G�&��P�/<�!>>O��H�	�����e��RH�.�/�$��ZҚ���~L1�{�]E@1�����oL��ӌ?F]��ԢOQB7\�b&���$h�]�M�\������2_[���q�ã{8��'f�q��b\5��7�ћ%��2Ð}���9B8�����.��M���z��%o��p����e�6�%7(KK��)�3��kr�ZD��]xZ���Z�+c��vk�b=�v|㴥.�MɁx��.;k�B�q?�4�m�Τ[#�Bk�-b��c���ۜL�&8B�pR�f8A����
�8T���$,�og{���@��C�<=�+�sp����o3%;9H#���K�u�*�KB�1�S��t������̏Ͳ�q�i�͈�|���������*Jy���MuTc��0JV�G�f�[��xG)�
{���"�ݰe>�Cf$��S�����Ǩ��t(Ѡ0�Kc�3����Q�ӓ�OW[r��g/���/��ޢU<��20۞1�������"ы1d,.�t?<��P��)˲rm��٢6���B���}bn�{����ŶIV���~��i�����w��~4ҟ�*�c�y('�~<L6u�MN�,� "�Iʽ� xY�sCWK'\ӨT���Su�8�Rk5�;1�ٰ�ur��������8�z<�kvn	פc4|<\WX"����%ɫ�KW����I0�ڑ�t6ąN���7�<�k�
�);y�\�R��2�z =��
bHa��� �$�������);$��w熓vK7.=F����Eb� ��MP�������tDy��V@?����O�Y S]>3:�Bt@̓^����C��k-����z����!p��	���vK��b��^��$D�Z���f�����X�Ho�L���l%��wk*k�pO���kY�M��k�����Ct�W��G0+8j -ƙo,Q�YߟO�������H�?���Sqy�eĬH>دr���u��
�׈}�nY�|;���	溟��$]-�� ,W�NrjJ$�ɨT��!�])�z?��U�i�w�.=���.���RE���+�7U�a�|�\]ѯ�_�w�n�p|V�@h�1	�ŠԠ���C(_�k�C������^��!g����$m\9��_��-񏈣a
����@��@l-l�N��J>OJ#�	�u���Bx��sTn#�Xa���w������U�O�a�lE���_`��Ob�����e�Aӷ�8S���s����y�4�=[���&h����M��W�L����g���Ok�K�=��y����^;�+�;ES�dIúh��� ��Dg�o\���g�<������9Dg� m���'���<i�����t%�X���o3��u��,�f����\�-o��������'4.dbUٓ������P���9k�m�W�xl���'�@	&�v��h��$υ"+��c#e��t����{��"3,;/5t�c�1��1	��3��s���.�k
Z޶�zW��!�X�) 7l���	;�XK({�g�=�#k��_��?	�qW���.D3��":�\(�h�Y|s<�7�	ܐ��쀹f#\�-w����j�gL!���GE#W�+�[?�g�q�Udg�bW���O� *a����1���f�#�9���-w���B���m���sk���6 ��-I.��n�?LR�3|��2��Dӻ��bɘ�������;!��ӛv4�B��1��U"^5PK�)"���Qv��܉K����S-���=���,�I�&˞o�9v-��U��i)�%��O�V%�H���ߵ!^�қ��𹩘��c�&��@��\��Jm�\(5s��]l��ǫ�`l�1f*�2��@�%����5�N[�A�E4��fHRq�r��s8 	��^6ɵ�1�� 0
9�)���G�L���^���n�?T�kW�a�y	�q�Q�X9�~$�D�v��=)_;�4¶9[	�킂|��c��"1��w�!ʖ���Ҡf#-B?����fa�4��~�x���ejY�Ac�rb?�u�v��$�p&���5��KJ��1$ܜ��l����rI�Z䝢a����۷f��M}A��s}�k��PcE�W�o8��9��i7��w&���@�ȭ�(���������Gyh�l���B�EL�T�"f������緄�;Z)X����I��֯ҽk*a��z����$��&��_�͕��9���<ȅI}q��%��Ȅ�Fw|`���m(�21{�I����>�ď��Rf����*;�(��ȐQ.��k��m��r�h��l/z��i�t㾥�� �^�*�cCR��r��eʘ�d�Y�~	=�Jƃm}�S+Q��aj& ��Ӝ ���k�*��ܹ��p�ٰ>�(���&�ʨ�l��\&mݲ^�2��f��P3T�uo&��]���dp���`�$�{������1twS(�,X_���=�����6]�W0lW�)H��PG���=��]���*�>�w3C9���� Hk���:�Դ��/;X�/���Cw
bo`���p�%�I^Q��g�mStg�s�P�>D|�v��i����^���$�|D�F�ܶ+t��K$�kl����F�2�R�/Ɲ�P�$F�P�S|�\�n��ע>)Fa~
������O��ˎS4;�b�[W�w2}��_2�0��5�B�Υ�M�Nt�X�%��= �t��13�x�`�n��3�&+��?%.��F��+��5�(�C�@$.��4���Z�������axP����?HOI� �B�X��ͬ���I`+�{�$<�	h���V��\�66r�X#
Ʀ�)ڶŹ���B 5�Ǐ$*� =@js^0���|��r�x	�n̏��b�D� p�/�+6��̏Bǝ%���n-"3arĻ��z�����,���ǜ���K�\�4v�S������e��M'Tt�?Uw����3B��5G��򦚇���\��٦wd��!�%D����K���V� �!0�����p߮ಽ�����d,�?Y��:��¬����Q��^��_�&h �'�ۖЫn��G=���3Lޞ�7Iu�s}q󢭺`	[y�f,�@?%�|PF�<�v�}C?H5�c%��'�L0�k����<�w��-��Ie�a�(�md�6�cH)��_�����}�^4������ʙ���S�TH:�dX�E$�!����ds��'$�6ԧ@�$߂B�;,d�)�m��Co�S�f�s���^[�1~����Z[gag��	��I�y�.EH�fKr�%��h���8D���43��!a\��lB����0��J8�8�����9SN�oCٺ������9�V��]�Yʲ�~My�E#�X�����ͧ��僧�w�h��M6畇 �T�!������p	%��s���QPT3���*Ȳ{�ւ�]A���9V�>8ڶ�]q��"�:G�#�uu���N�'1%��[t�~]���7�Ef �Ⱥ[(�o�I�O�0��p���@��}��JT=�|�����h�hr�n�.��Z�{��C���Ѣ��џ��BE�g�ܤ��/�t�˲@�Z����O�{���b��\wB�o����ʪh|�1(^��A��@N�i�m� i)w�1�ݴD������� �e|;�ی�J&"k̢^���UBC�]|#��hJ���9E��'ƞ=\w��X�ʔV�
�I�yQ`��>�@0��^�i/��ً�yDG�?�7�mr䅀�
p��&6p�ܮmѼ+����z��<.a�j{li��@s/#_��ϼA�Nv�o/u:uLa�*�/ս6��"~ee����mț�i��i,�"IUyk��C�E�XHŠqh��D����T/��b؀h��&�h�M�&����y&�#��6y)F��I�@�Ŝ{��U�aB�H̐'n�@�7s�B>E-E^ڃ~M��=����_Cu*L1<�?� Khj�,�M/&���}�'ǨU3В9�6��'G Kt��e�V>�+��0M��* ��|&~�Ŋ���k4ПäR��)HB�|�$j�/MƖ��3�]oK����Xu����N�T��A뎠J��Ľ�e:���5��6I$��1�}ӵ$KA�XT(ܬp�aRxBc�?QO��g��0C�z��U���̷$S�!�袨�Bb�l��ɻ�Lj�$�"Z�@Π�|쬬���<�ѝ>�Бv�Ĉ����
�6Pq�pN�=�sSZ�xX�'$��}As��^��ҿ*���衰���ȗ=�v���L�����J��V���7��	�Z����~p�`��P��L/;�kǏ�����$$����H92� �A6�_����\��t|
)��pf�G ~�~�mȠ�$�T�s�+�1{�L�^�J%� eT�q�d��낥K����^(kb��g>"鎱�������ʋ������	T�-�nC3��	-�mA�ΊʏE hW}�?�n���%������	_xz%��v3b����ʷcC]�u��#,|0�Un����$�ma�.�.Pk�NqA�����U����49��ՋA�� )k�TA��q͂�
��@����g ����WM3�Ϭ��´�ct��N�x�~� �q"�.�'�Wo�-��	�U u@ts�����ʏ������I�,����~|?|JKlH��t��?��7@&��J+�ֳ>�����)�M8���j5 K�\�ϯ����1hg�����@�	����S�)ܩ��U��̒]	����A����6��6ʲ:�����3};;����+�0N��R!'H���>���w�����:�
����9�:t�:M�C��T�� ���er�yXB���k?�]1��ރ�6[H1Bx��Ǭ婎�Ʈ�+���O�F��UC��
��o�6�����O����=�iwE����){�=G~{�kq����#@���Ys �*b@��L�%�43���R��}Jw�A6��X��0O2��Hd����X.N�Y�i�@�I��l�,0�s���U���ĥ�������|����1�r���j����h��2Rرa	�i&cG��mh���Ζ7�4%{+	5���!�=���d!G-�Xy~���X��l�T�~4nw��̧�8 Y;��	�2�O��<7<�ψ.�*M%?����-K��d��^�\i`&$/�/aV��JQ�Ӂ�U�%q���U�o
��1��x 0 ����-�/"�ᮊ9qu0>���A�__}�P_��ܘ����/.c��k�&JSIfDdV�έ�bR6�#UR�;q���p�lNsι������ ɖ����U݉� fb�Ç\E3��v}��$���B٩�b·��|�C��
 ���΍Uc�!&I�J6� 5�_4��w�UQ3�[�H��RnƮ������%^]�N�$���@^}"�����e�� ��6��N+u������	i ��J���m��4����Z�}�p����B�sg ��&�.�`��`�r*��X���
�(�y�\k��F{3%iֱ�*�Waj2���z��$�d{�0y��'g�Zp�1�Z�\۝1�l�ܭ��'���v�r����[�1��(D.x�O���rI8�[���!��	�� $�mIg� Ҋ����>�LT݄D�?��sS-55É��b�,��1�캡���Ao���!Y�0W��P�M�)���9�V�ׯ��*�m��h��*3S0��Q��jL�p[�}�X<�=\v ���-Dُ���i|sDs�%��{��w��r9�j���T���^ޙ��T�����D�Ҥ������{M^|�������������Z�	RVz�$J۷r��$ɏ`�g3�����0�zH�>괰R��kg[0xr�}㣑�s���a�b���p]:H�O���6��o��t���cA�$.(��I�Q���2x�� 8�O��i��Z�Ŕ�Pg��R���.���E�#�Z��8I�E+)�4���]U��S��A۳\�����Kl`�E��b���J�ѿ�F���4L}$"����I\� ��S9/�t��T��Y���Z�쌞d�1�����O���v6Qp��s�ִk�Z�b]��V�N���,M��]9�#���(�[��OsP���Jt��$C�GK�����(�k!��!DO�<�7F*��5��l��tD9���l���BN�V>n��
^�ã�X~����탑rˊ���U���R�,�8�'c�qw4���v��A���]�hɯs��/��:����	�"�`�;,~B-���<��j�AK:&�)'0��;K����u���
YZ���Ņ�u���HSv; ���������� ?�ʔ��F���dir��ᅁO��姑��C���CY�)�j|�N
�"m��yɎ'01 簒q��S�\2#&��&1(�!����s�Um�Y���} �?��
y�NF�1�%Q{�B���n�*����-q�.�<u -�_����Cl�~���$�!P��M�l����v�z�8F�al�D�`�'l�����b�,�hcu%ޮA�?��DA�6ՠ�_��Y�`ӈ�����U�O��h����C$v�#'2���\6+�SFَ��V1A�k/�#�m00�6���B�]�f[���kH��绎2�2H ��k�3��˳�I1P�(�i�ٶ�͛K�c��b���c�爛�>�-�s�UjCS� �;���F(�5�5�Zm���l^������|J��H�r��	����vp�C��������vW�F�����B��w���@>Vv��y���]I�����KT�ڇ���"�������i�ą����d��
R�ŗ�4>���7n[x��j�'T���ǿ�#�Bx^-�3��=@��3���r�Xz�4)i�2�yY�:f!w3HS��$Ӊ��b�S	��m�zcMI qZ�q`i5����'\w� f]�?I����|��Xm��������6��'J�_<��5�D  �Ȋ� ����<���I�3�4��~CeĴ�18r�m��s���p���n�ϼ��Ѿ�}?���YA��^+R�QXH�;mly��@�:]Ҩ�I�/�t�.�sx�ҷo��t�YS;�f����w�ӛ����#qO�m�_\;+6	r� �.������qe'w|�`�)�B������Ų�'w�ģ�xUk;�k��i�'�A�����v|I��$4O�ۑ����D��(�N�k_��T`rH��V>���(��ql�Oi
�������{S���d�#�t��X��}�V�Tt;�ݘ��Z���I������d2iNs�I4���N�V�������Zpw�w���N�&F��Բ��R��O/i��B�i��=��?8C�Xf�mݏX:��[�wh�ϖh���4)定č�r�(4��|JTX�9c���;A
D0 g=k];���]%l�#g�4U�O�f��*�}۶���E�5���Y
�OH2��H>�Zr(q5�v}��ϡ��V�Ӛ��͕-��f
ݰv�BNN�hѺJđ�p�2)�&���S`�'��s`C� �kI�N�����f<K4��c�Uҡx�#�z�0v�'�9�jŧ?�c�E{3�ΩgH}���A�����xL�f��-�zͼ.V���j�j_�,�G�׉�A墨P�W˖�/ڍ��w��@"��~1h�m�#Y|p������ܿ{la�%�b��t���`�g�a����-?jǗ�o���BCu����r}�����y�C�q�@�9�H��;)���Ϊ�����3A�Gz~>uώ\S��0����T��_��d:f����y�Fi�:���Ǘ{�0xz�׋�R/s�OvrG��i��Ӊ�Ku�����8/E+D���'f�_r;�~<��T-��>�+�s-S���%�������`�ٳ=��8�U;E
�<�c�ru���YA� 89�9*D���ˢf�V�et�>¶M�� =v�q�%j\�c�_��Xj��Ǘ湨ВH����<�B�e�fM���� ?�B�5GI�-�t��IJ���6z�����f^�����L����B�&��(�D��P��*����dO�H��(��p;y�ɽ�҄�VXv�x-=���c
���^�t�s�}�$4sh�!��!�' E@�ؽ| $�y��M�+��6g	N����0�w*��a��n�"�Qܷv[v�<Vc:�"c
nA�O���B~�W�i��Mz��ݏ�k�Rt�����)U|J����Y]vϋ���B�U�حl�1庪���̩�e<UV�ү!�ܮ�F`�����6��.4��0A�9�x۠1Bol���ĺ��[1���F�U�+X&��9�i^��/4��r�VJ��c���ݴ�|�k}0"���{�亨IPwq��!u	�B� ;�!�V t�J�Ĺ�V�]��?iy?�p�R��!���z�*�d>%��=��Z��e���"�Cʭb��p..�X�ʿ���}Ta��K*|�O� <�Wӂ5�(����Z]�Cy#�㿆��
�Ғ�Mm��X\,J!��r�I~�6tr: ��珇f����<-/�j�<��0�)�#r��ٲAZ�$x~3]�>Nٖ0�R��@���~ɾA�$� ��wK9��jB��x 0���\+?�йޮ���+�g��]z�]��n���np��2��6��V�E�^�ڼZ�H��{���������gۥ��R�N�߁�	
r��}��O+F@(`�ɬ��⪙�-�x���J�Ձ�f�Z����c��$Lԉ����g��Ld����V�I>@�S��m2t�
~ƥ�z�Y1e��$�V�2m��{�ŵc�1{h��{�ȋ�E�:�%��J��W�� �@� �8*b6]��"��S�N��_,���r, ��j{�N��1����Ź
�IE���P�Қ}�ii�������҄q��!|u�"��X��6���P�AkO��.v�{�����[�uT�5��P�H��cՐ�`��G��s{M?��{M�=$n߭�=��̬�����
:&g>��E7)'(�Y^nڝl�U�6Ib	<2�d��v���yZH>N���DCy��&Ku�z�����#�`0�D�m��+^����:S�� 0����>��v<�>�/A=6%0��OErn������I�"�\�HŰo����Lvb�d�^ho�Ͽe�E���T^�giS^L.�#ؠ���u�Sr���i�cy$V�椮���^ȿnv)Pv�W ���sl̾���m��+���7;"o� 'e��yb�B�m��8F1�Ԛ��ԟ���O.�����~|}R�p8����VS��
�X��&�;
�5��qs��i�!�!王{IܐB�4�:�+o��
�֯�o
�2 �`���}�Q\͹oVO��9�縺�s���H�FR�2��t�2D�7�p"�ۮ�9�n���C��c�.F@����+�(��q�R3�SoK@��H��\��F�(i5�vO�M�K-�
�����~����bxxD�X��<��jXk�M�����¹� q>ʺ͌B�X	3M�u^nG�Gȡۊpu��lVR�_=5���&O2���y�s,�`�8В�,
�ˇ��g�{N|�E�G}[&Q�D<px�ruN��{bѡ�l �,<4S��N %�J�t��lo�HP�rc� �\��\_+��I��)nY��|��r�%�V�*��Zޢ���eQ�U�Z�I�n����L��J�)������lpX�O��[�疻tZ�̜�]�Mv�7��"I������y?Hmr�`�Rye�	276��%���T�h�꫼e������~����������_�����������s�&l�����Ԧb[����N��N��H�0<#ˋ��z�4zWA�q���vp�0�T����,sYG*�ߛ�+ެ�D~�x�t���������I�ߦ^�,�>�K1� ���z�����ܓơkf�ͮ54��@��f����6�WL��:�/�}�A��k��]qOrq��:힜hn�M��l����e��Z'��!����1�]����c�*����n�u�W�O봣)<y�S33z�C袑�����.C`�Bam��|I�=O�����͠c�,tU��ْ�NJ��o��|�⤉���y$ee�4�e�/�E��k�g'���_\ﭬ\�)���~�z�K����u�j��&ƿ�FG(~�H*昃��N����H�k��l�2��������`��zd�T'j̥BNw��6$gmB[�du�j֛�~�DL�O����5F��覸a\ވ��ڨאqEy"c�j�K����
��j���>�6�}��"u>Q$uU���K�Ó���ϑ�\Y��������9:ecd�`����
�����D� ���(�2��1ҝQ��=E�!I�S����/��)[_�q�hI�H���P|��X c2f�qb�su���c�i�a��!��'�@��=�l����R�蠌�Gs�������H�c�хN�85[�1�N�`ry�����]�^:�u�����?Eu(t��ч�T{5!�-u�)A��c'(�u��U���c�n~tG��A(�=���_ە~���0k��3 �g���^�e�>4'VOM|�ӄ�'B��K�}/�%�y�+���X#Ջ��dK�D��j�9h�V��UG)�&�չn�����*ra`
5��n�	h������G&
<3��3�s:�� VH����b&X!b�|��'��:@�z����fQ���P昫65��}�˓�{pW��8$7��uR��G��]*��K��KU�q�|g��)��Y�k�xa�'P��G�۔���eb�����t>ֲɇ�Es6�V�_(W�Atfş�����z�5Y��߭1V/t5e.��+ h���[���7ܨ�#W���N�����w�]
$��(���?����0˦�'^�$3 p����@�q��$Ƨ��X"����-���N	A�Bؠ��L"����n��E��S�����!l��9p)ƘC|�����K���|ȼ)�P̩-`��`Oy*�!l�\�G�􇹟�!! �W5F)Ǟ�[���mi�����),h���Gy>.3zx�tQ�:P�>>3��W-�c1���&��ԛ��sw'Pj���ԧ	�S�Y���Æ&]�����CI���B�P�L���q |4�p�e<LP6����4ܚhVH�����h� �	����
��q㶂ƙo���ѫ~�r��ٳ��j�.ă2�<������^w����?<�1?钠�P;m�<�W�\�X&�;��\�F�זoo� k<]/^L;�@m0�c��M�7(������VvIRF����ц�����!����i��qb�s���ޠ���]��K��h=T��7��A$r�5�����ӥ'�L���/�KN������c��v#]2��?�gt����قO�g�=˸��ҹC%B����!B)A�lW6��|ٖ�ոA�%r�TY��f��Lzi�I4����J>Fw9����K��Ի���*�{�|t.a���8.�㵀���B>�h��^�e@��%u�"�N����lqPLyP�������Gf��B�{h�ޡ��z�3LM����*�ڇ�%e�`7��G=�Eg�cl���v%�J������#=���&��'x1���{��~�@��-z��x��8���(8s$)��9�?>8t˰bv�����,PR�A���p���$�R�����lC&ec[t�N�'^�<�-D�^�!X.@A�Tz� ��$7�8��z����O2ϯx�D+���r�&0mn�I���ӱ�*��A1s`��뫥�E4�{Ax�tXT���;�}:���6,�z5�O_H�_)�lF��u����̂�&��ـ�������O����|*��-�{�x�	��r^����O��T+���K�)%�������׍7��<l"1�i��LO(?��UC-ٗ7�w���UԶ�)���*&e �V؟Dh���v8�J7�t���k:l����"�^�û������_
Ks�鑤e���<�u���M��L"���G{_+Z�:������1��?̿<���j)�2��^�a�$�08�Yr�<X3�=औw)�j�9�pqm.{_�O�L�i��lP%L�Sw��b?61�E� �����e�f��blxb�_�M\�)�~\3#YC�ĳ��D���)$�<����Z���-��[�[2�j
�0�"H2����&�����{;S���?%�!�*���=,��t3�l������w�m\���n�i��n8�n�c|��mù\H/���B�I%�	���k M��cى��F{��v��^v�-�+������0��v�����gO�c��if<�Ǹܓ��C�^ v�o�8m��H��i^�#-L�Z��ߞ}���	!��i^��|,�7!��ȃU�x�z4��67�O�f�@QQW��5 ڮ�%+/3
h�[įj�ŕ�`�T�ή)�7k� ϫs��LA|O(����|�\g�\k���2�����ZM޹:X�)�Dq�0ƟƜa�dN���*@;���1��@��kV˦R�qv��B�������+Xݫ�[�G�{�b�z��i(/d��!^Y����9d�:P`��d�\��֨�q��4V�s͕�$US�x�ʘ�:�
|�ɒ���b� � ���Ѕ�c�D]L��S�0c���Y��� �m,A�9"x��y�J<�y?I��	~�W%B�"�7 �T�ʮ��ե��k،l5X�`��<�\d��7��nλ��kt��#����W8�8�ԉ�{*^z�J'@׀� aJ����_���9�;D�Aּ����>/ⰆD̓ǎG|K�tCUƵ2t��xH����s8��6a�<?����Gh�IVv1�~��'{�dc��&�*Wڰ���3dKB4;�g@6'�G|�X3]���*���F[�c]9k>D�U%U��T*���x�xBtFNޕN�BA�.+LQ�];�P�~���d͕F�hۓ���\,��n��*�ȫ�V���zs�j�Xޘhz�n��gk�ևE!6t'����ڋ�����s���Y��-��A�_��8��Jc�ld-K�v��q=�+���;��|6�)�y`7��rM�?�-5J[¡˂��ONEkdu�ޯr����'%�w��p��8��p�C�����Ҥ@�P(�j�ˑ�E��r��J]{����&��A;pn��g� 1�
��[�&ؠ���j\^�Gb�y�s�N��|��Hݼ�y����<����ס���FLl"Pltb�f�X���(��f��gsY6��T]�̎VmH�y�W0�D�4��eiY������j�5%��y��ge��J%��ݬO�=}��#���K�3ET��<+'A��%݌�2��lo ��U�2�X9�ٓMssW�Jk]���|�)�Ơ� ^�\�e���}O�1q<����r2׍�y��4�Ԛ-��.M�(�x�=�]5��&A��o���]y�O]�#�������4$��|������V�\��Ԍ�����o�i��fMRkz�F=.��K��p�kx����Xu#��҅ 1�J���4��}
(��(c5��;&��L�:3�+mE�ѿp��_�{W��WMy��9y��(�ҥ#��J�х��@��m}���fm^��{?��YKGc�.j�=J ���In��A�{!D��_�T���H��G��v�6������A�nuǋ������E�+�{�#�)y�S��nnȚ�Je���.���Q��kBWN�����8��=vY&f���[!�GA"e���^9�l����'������F�o�|�h������Aԉs�W�8>��N���{��uKW�s�p'R�Ou%� �Yݣ)"3H��S;���p`S��%�K����k~�!W�������r��ݤM�C�L�SE��"����E�����\6r�M]I�f"�%H���Og4��R[Hk�qqq]��c9�Kh��S�`�PU�^�+����sLϻ���|ܗ��w̒���% {R���He���#e ]�Pu�˼���ըgI+|�����]_7���j�Y�d]K��+:<c�q�1܅c�)�7�,�h��x�~��d�����M��^v��c�������6W�*B���٪f��'�;�q S�y�*b\�|"z�.��ܳ&N�p������W���<+4�1��T'SL��?(W���c�$��a�Q(��A�*
��G������Ƽ����ḧu
�9���|e΅G�aq ��3w�"3qԇࡠ�|M^��䥒.�����>�]���07�ɜe�3�}~�k���D�O��C�=�r�'�����L�/�q~`�C^���[����q�ǝF(��G9���r�»�6=-�0n����Y�lCõ�,*A��6�9�X��'�ޥ�E�T�c��R�.��!��00-)9�����7�����{�	��0��]�!������yw�_�������t�.9N��2^���P��{��F�����ȕ��+@��eq]���ĩ�� `�����]=\�������<��0�l����f@� t�g�oyן�2�a,��U1y�\Ԏ�R���G+i���wݼT{� �lU���k
=�V��ug;C�O�X����q��[������^(K�rKn��c���͔�eK@]�s R� ��"�+�#�=f���Js�"GC#+#zd�N�4��^8��G�&�*w#�*P�ZЪ'����F�m�F������|vؚ����#I�Ԓ�|�H�'�{5���ֺ+SY��\�LHQp�����
+�s,�FtX����.��C恼Cg4ĺu�~��k�� @���x��`ڃKV��FpXZ���O^C_Y�٥�q����� s�ی/��{��� �;���p��� ����m>er�N�)��C�j�BM ���qY��|�����q�YG����Iֻ�3�y�In�äx�e1s�����~������M���2��NTM� ��2�O���S��J�캋��u�X�/�^Q��ں���Y�d����{Y�2,����w��#���*�HV;�J�71"c�&�x{���q�Ѱ�r�&30��|3fƷ4\��r�I��O�����S�C	��}�!:�Q)���ZZ@��JV1xi8/'s��ӿZZD_~���j�'������w��j:�Ĵ���Ä���x1�a9k���۲��*��G�x�4��8����$F6�n�F -b�)f-����C���M kr$�G��������X��t�JH��6���!2O/B��>A���E���b5	�a9B�M
� ��Y�ċY�0M����c������t��tk*<����K�u��2�!ɚ��2��9�d��P�+�\����%�ol%i5���lZo��? ��9"\ �6Z���\���F�)�O�G�+8�`"{^y�
��c�ݏ�P	�yu?�s�	����RAj���7~ٚ&�'�,���r����)�fW�=Ք�����z	��ߛ��J�ǒ��C�S��VE�h�ᤞ��T�.��XEA�v�i�� �9�!2��%&?m��.���I�m$�v����锈C��Fp�8�
� ��y��H�8�b��w�����O�	�Z��RMpf�$�	z!n1BT�d;d�ә1b_���S��r�)����0ۙ�Y<�PFb�ER���Ma����B��pnR`�/��E�1�֪���NL�`mlpM��&�5Y �~AH�����J���GL���꜄LD�j�uo"ul�>�f#`�(6־����x?vۡ��ޜBb(��x�t	~�_��Q�S�d�`�P���>���ߣ~A�+�Ș,pJ
�.=-�a�m��Z���qRB&gB��I� ��� ֑�x�G�Uz\��S;�F�h>��B�ĉ��p��u��~�"�eu�i�9�M[�=��{�$��ګg��	��9���:'��oeI��3�J�"�s� ����W0�K�������P���@���c�Nt>ѻ{vV6=p�Deh�P,���͆`N��uj$/xcO��d���[�1��H�2fc��,��}ep"���ʤ�#F�p 3�H��y�/�b6��S�?��7�6[
u������{���qx-�`P�}z3�ǹ� ]�!�ݬ��ˋ��T�!|�E�]R�%tX�m���97C��+��ɾ��_�td�p�t��Pj��,`�X�>�o ��~��+�!�?ItA+�Zl�v���T_�qŴ���~q\���G�����	� F�E'�³��+�
1:���z�k��E3;�g8��3qh��� ������'g��*����/�Wl��z��鿹���Θ�-۵�En�&B��� ���4]�����<��K��e��K��DI�>b�<��+|�S3��7��᫑���y���}dV���0�^z9��<�u��[cv!�p⯚ۻg��������SC<�h<��q	�����JKvl�ZI�V��+eVQ��r�6��q)�\*����^}b�5�X�nb�8�n&�5��=�� �G�A�����nC�Ygf%��mLp��%�7����n"Ƿ���Ww̸���Qa*���~[��y|!k��p
���e�Q��D�ت�z�6ͥΝGu�[�*��`_�,*d�tJW,�@rߎ���}8�����w�y�"�:��F8��Z8��ۈ�/�O�AB��,�έ�W��<�F��U��H�N�F./�8����6��tVf�瞣u�4���i���<�j�H��l.��=�Oy1���eV�<VZ�����\�����nJe���h¸Nl�&9jvo-W7��_	,_�2��'�ǡ�if��ݬ:���=����B^�_�5t��R���#$G+
������^�}H89�"���	-�����s3K��U�V�t�@)w�z�v�z=���*��<rB�V&���K b a�԰���)��Ȝex�!i�g�\��JH�]`��(�J�%v��Z�VH|�fx"Y�ݣ(mҒs�H~a�ƌ�C&~������dP#P��U�$�Q��Ǿ}԰�`�$�1J�j��k���ߑ�JU-�ivS����xtKnqx�f�Q��Z�N+����q3��d����(�[�j���~��Ҍ�B��Q��sL���w'o�#��z���
�tt.X�2�����\��?ׯ�[@�$8�I�3]������ԩ�H3�?���!����0z��F��VQ�@�#����&$�9qL���ۅ��q�c���(�i`�P�!z��+Jm�u��s���n�j�j��A�܀���8նn������0!
`��r���N����*�Wv琵� �����vqyp�u��c��(�ӊ��\/��_u�!o�/��N �ʨ;��
�������q��E��b��Ͷ�r_T18��v�h��!X��\ʌ�q¾3����S���h=L�����.�=���!������ˎ}rVac�CW��'B��]O\�;r�/��27�S��ʩn �T�xA��-f������Jg���L�S>��Pv�:O>�s[�
V�i�6�V�,��+�5���o+&���Q� ��%����nR�V;an<�#]�wN�Η�2n���?������z��H��%·�>�`�`y��1ʥ����AmE��`�5���/8��HJH�F��q[�<`6U8{���t5�M[�#��$��ц7l{��ןi����d�,�5�2ؼ.* H��&e���y��_�]�O�Ԏ��70�ȷ[���ߴe5čP[�>�%9O��I��B������؅�N
������/��b,�ð־��->���(���%ت	�������}��

��}~P5(��
E܃Na��k�V�E�����\D��/:��2j�sO\e��P���f�<4Pz��x�o��fϬ  ���Y+`W����I��KEu0H�uXb�V�z���-V�J���JE�-nO*3����n+�dF7&l��?,H��4,�U�;	)��>i�q(�@�7+]����80ʹ����H�O��A��m��{�J����� �:�A�^,�u�'�����|>2�rp:��. ��Lt=p���E��[�_���٥�3 r\��+A��@i~�}TZ��l�.����y����Ha�M�4�����L;^�>��C��΍��P�8Su�6<�ŪI<G�Z.�i_M�39�4)��B�T㶔%��U=:/b9~Bf�-�h����_�(8(���w�Z���
� �+�o�,���2_�;-��A</p�jl�
QBa����Kd��X���h[�����k��q��ɋdy�[)H�:��v&r�vy�ѣ̚%�qk���)�a!v2Bm�)����%�κ1TJ��hm���x��@�CWIRclϓ��w�YHQC����x g��L����A����F�C+�u=��,WfP^��d2v����l�g/�L:L-��U0q���$M:���"5HZ���,.hK��Y>���L�����LI�'	�����R�ݫ�4�M��/���iZ*�%܂�_�ŬCK��W�(�&�ʠ�|߅��I�p�'�kz�<G�o{'��h眤s��<@��;���$�( �񠹞��� �<oԅ0�U����#����5s0��������#$Xc-7��y�Vh����u�x��m��S͒mz�q�j�&IK3ʧ �Sd��v�d��Q����v&�Nl6G�w[�%���X8Ut��=�ܐ%��Bq (�M�YK��"��C �&��Z_زM���EsbIK
:y���a�����;&�7��^B9f�����V��Y06����;/y�k�R����ߦ;TO;�,FCu�f4\F3j?i ����^�jZ�z=�B�i�'��R�d6���Ϧx�w�q
��۞yV��@`ye��E�M�Ҭ5�q����A ����:{E��,We\��nґ��y|C-�TՈ��� \�(^}�^}i'-��b��'��Xr�)⏌E�9���9�����w��lJB+x��W�0�be��4r�铠�������D�ƻ��fx��H��b���t��L���/���Ż�0��pB��g�ֹ(d y_��KR�leV�wᶅ�޲Er�@��u�u@���)��=M(?po����sv�����5�Ε�(�D�q���>\�߆O$k&SHD�Bzd9+���+�>�۫��>��gH�4��?aL]K�T����~	�����	��Xl�'SN���\�<�ϵ�T��5�r��)~Ć_�A�Z!�����>x�������<�͈�+�g�|֚6�������G�sv�,��-Xxz�B�N4�+��@��}|�}�T�7?hǉ���#�����2�_�)��l��|�&��M����I�k�_�u�|�FUt�Z��$P�*�Ȕ:)5��N}��Ͻ��]�)��)�box$�"��ڋ�K�x<�S�������s���v
�,�Ak�6m�f���ey�z=#/���{�':���t�^ݘ���c쒖�
HT\�2��
N�~����Q����*��B*�5�읐r���l��e�"8�X+{��P�da���Vy��%|ʠMg���7qh���}��M���~�p��S�J[;ۻ<T1�j�9��Jш����DNC	�G�r���t�m4�����p`�fk\G����Kt��t�����.����\?�����Ml�����y�2sK1�S�݃-0�7B��ma�E"'�p�7^aǕ3[���C��8��B�2wɜ"ј�-;���'����3��Վ��*t֭(��������ݪ���w:�?H#ήj>S�o�'
�r���:"W��9F���V��Hl\�q�pS� ~�a���S;ֶ����p�B$2%�K��k�G�`��G��3	�uҢ��l�Ԯ�ָ��	Z���`I���ܽhh�%ނ�ܭ	$�xNo������K����U��浰�r��K�r1W��oI/�������H�&��n�joѲ��X����" ;�	Y���m4n��3��A�+�����VSP�mE{T>4Cq��<&]�
[�|�܇-�ٶ���G�(���n�<?Ј�ϘM�B������[�.���l�;(��p���A�s\�R⑵����rgk-��K�����|�X�$�V&�����롴9ov�����T�|� ���P�*PK�����m��<��-Z_����i� ����1�c6�dT�P�k�be�Xi��~/!QU�d��c2 ���Lm"6
������g�\s"�Uv�ڊ�ʧHԈ�Hw�?�m��[n��Η��\}qC��:5�v�R�W�~��\S����J�N\�V ųHM�$���1ML4�kY��x�4�<	O��2Ň�Lk$d$�̟}����<
����Z���wy��9}}�Zʛ/~�f	��sB��m�t�� �g���t���<��C�{���a_B)���и,W��_���G�l�w�� ��i�T{D�{��}��6V�)�<���ZujT���q�6�I���RZ����La(���'�<��=�Z;E��y�/��h=Y�_��y:{�! d�;�۲*��{��)�f�Y��T�:���/$	�Ȗfi�g���}�<Y���[�R�m�x��ss��z����D�MϹ�]�o��ےG9*Ȭ��@��
Z~�}�(r�/c�OpE�@;&Km�9%�b5���J� X���m��QW��cO�+4��ƶ��Z�������!�U�M���C�I��L������Ŋ7�SOÒ�.d Q�KcϮ�?���/���qHIa�k��	��+��=��;z��o� ®<O�f��e;}/H����E�j�����T��Inҍt����<+�z��Zs�oE��(��=&gvP^�7�oL މi��ǵK+T�^'���z��X|gS��n+2�I�n}G����	Q���P�~2��8شQu��J���B�C�@��EO҉�N��
Uu_y�߱�Td��7�U
|}5f�+D��<!HO����i�@f)�+�;���b�n����+��,'�
,>�Z������Q��k��t��_�"���G U%�g���eJ���4._�
ԥ�����!�\H��%c����<0K���m�I�CO�,�S��W�]ޝ�ބ�T�LzJxhl�-�~��G0̜e�$�G�5�����^c�(�%x��0�S�0��ݖs>�:��~�{�_ˀ��2�٬�KK� ��F�;:�.N�z8ͫ��W�{�s��@V1^s_�e:G~�K�Y��i�t	K8!����Y�C��=a��%=|��ˢј�S�ub�:��w��n�0̘��(�0"m}2��{p����C����s�8�� 
 ��-?�ᆧ�*gI�R���#^b��19ĥ��@Q�>�V�8��xBy��A�X��=���w�:�'F�k�ݦ��ġ(���{P�D�\g/�M��`JǞ{�s�Jk��&��d��P��J-w������^=<�*���*�_#N&�YX@p8�S\߉�����5�$lE@t��Z�f�I'e�k�#��F#��'b�V�) _��Y��n��e�� ĕ2���>p�{5�ܪ� b��[2����2�Z�?S���g�X>D�X�=:�����tOJql|����6"�S2:�fj�|݌��X!��KP���+Emr�%<�gR�������l��]k�2�dF���?\!g��A8w���X���nA9��D�Ϸ�����c���Xa�s9o��\��]�?�2��ÍG�+�K�A+ڧ݁"]�E��`��{+��n�`���M�u��!0�w��U�0W���?O�B��c��E,�F�7�e{8��ے�Ӕ>an�o�f�&�c��1p�l�ݜ����� ���c/A�SeWP�4x��[���X�p~�e�+ms5K�+���;�����=�'���`�Qˏ:5@2�?|��|� ���G�b\��;"��s�#���1߭��ͧ��$���o��%��5�Dc��0���&��S�M3j9)�kE���p���Ƿ%���/�QL~����k1��Rx%�[����y>��h(�$b�\Ą���	ѽ�qr{O	�����5-��QP�`�*����r�P�c���ۑ�9S�'��#%%�V߻�V�H��P��h������ʗ��"P9���P{; 3Ԩ����BE�]��l�,��|��CA������T�c���N�;qZ���n*��ǂMk��>J��5.��\O3��T@��\.�����#h%\8{�@,�vC�+��]����j!�q�� qǌA^t/�� E�}�n��E8&g9t�*������Ɔ��"����Gz'� ����@�1$6��F`��|~"8�J�x�>=]`�������:��}�(�A���Ǘ��{�.,й��y�7	�+.�^4�Y�u=_�>�k�D׼w�s\���8���D�;k#.��<�������=���9\��`�x�yG����b��5��CB_D�7���*ԥ�PRI�|^1���)�
t��Զ0���d����jw��(2�MlC7!� ����8jy(��i�	? _��Z�����Y��ǥ��!P�Pf�+4	�4���&�ό��a�b���­�E��=̉텋X��ʟ�p���W�Y¿���3�cPxHڰ��=�0� ���TSZԮ�W^�k�uN$L�>f nBdޅ��Eh-�+�����=��,��E�)W��̞W)c���ðFR��_\K�!w����r|)���2'�r�{����X-����l�y!~J%�`��jf� �t/ޕ��m��`}>-ٷ�4���t�Giт���I)���ٰ#�S*g��L<�WI��Z4�+�Ee�;�."t�O`�'{���3au������"��)������K{PR�Eа%Sw8�D�
�O`��@��iݼ�*�9������.��,���+�*�||)l��]���8t�kc25<�_
����r�!�_�3�/�P�q�9�m�]��׈j
��`�hb�1@�x�r!R0�}�gs��7p� �F���~*��0L��yQz� H��C����3/�?��O�� K/��OA��6���������.�Gm�!��N_5z$�q�ڪ����E��BM�1.#Qy�q��1�ԋ��1����"/�ّLQ���'O���
�����)���i4&IL�ANN�J����
�L	( >�/�4�Fe��E�c�+�ɓlg�
*y9r����cҒ�4Pg�4����UȬvʥ��@�=�J��쵵�Z�sT�%�/"��2}+Ek�o��E��Z��F^�$��iVف����3�Oy��J��@E���s�-���ˎ����U��Q�ӏml0
�)��7I������%�k�=Xҭ���#	�I+�JK�Lnx�
�er��Otf�BCd��/����-
;n��NU�h��W��Cc�W���Tä�»�����ֈ��5�t�Kc8
������;�?�^S�Rѩw��La�?�����U���X���G��#ǼO���j�>���:W�;�y+���c�3n)y��- v^�/!��.�q�X����z��͢��8Q$Mq���qu)���]u|��!R���p�Ut�i8
J��U'���\���T�D(��p;�t���Cc�j�����MH�-��FF���&D�Pd��tKJA6T%���z��(��:q�}���?�O2�;ۗR�AM������8wß�ńb�����&���z޻�fT���9a
��g�Lyn�DO��k?.S��6z\�.���'��������pJ��=�n������TGB4R��`�	���?�����c��ѩ�諒Eȍ�\���>�)Xj�	�ōCִ��hÅڊ�>c����� d�ԃCr�6fjZި÷&����6.%aF3��1��oӞ*���n����zM2MN�r4S����>�(t.D�8*�_܎��<��1
�L��FC�h:Л�4H
��ьd�A�<tz�y;�t�ɯs)$�@'�Q�������&#������w�l�Ha��J�N�|���<��/@"jv0�z��M,�c�#�8|w��mmm����Q׏T�׆�5dӸ�H���e[�H>�̜�^��/��0�I��PiQ^fP����p\��a������ӼDh��(�s=X	�+v%5��!��PM��ѱ\���j-�2Ǽ���������&�~�/˓�o��8!����.�?�Q�����B�����~D*IRNȴ��B�W�n҇�)Hm�	�`�HY�F#ȿrGN��[�m/�Q/4�4	r@\é��uO�(O�5�Q<��\���=��x���ڸ�քS��P���v/ݫ	5��J�I�OS�M���#G]�)%D`LǑHe��j��r1��՜�>���Y�7ԢD-�K@��9nAm�V������i�4U�F�Lꝍ���aga0Ћ����l����T�\�T��W۰��!Ї��ma}#tu�����}aݐ��,����{6�����[X-���*h��vo�	�k��������:�2 J��/m=i�[�I�G�+�Q%ަg�s��O�14�؝$�Kۓ��~$�O}&
�zT��cK�+P�$R}C�&�G� T.��a=�)��~�
 uD	f>��	;���̭Ǆ�BaB��;���W��➔OK�i���jɴn�-mY���ǀ���5��P�`����/Hl�S�di�o߽!���"���G!��`��v�*ޜ���ɫ�Ơ�g�h�'�px�
N��;�+��m �-��4/��"P	}Y>�ERb��^�aV�'X�R `_����U�����x�2��C<�qO��\k���+>��:�Y�_w0H��Sg�������C��7����5+�;�>���������W�L�<���5'�{��J�"lr�s�������ʃR�����4! �	���3�	�7qP�\$iv��fN\��Z�����%7��1��Z��
��e���q�s���5S���B
�ێ�����ݚ��n�c��fBG�Ό��E%e���F�\#��7�z$^�EC��o�*n��T�ӜD�7y�'t��K�|#8����q�d���G�x�I�f�Q��g�_톼?Ԯ���J���D0�k�n����ȋg$#`د�gQ��"��m��m��C��.���j画,����H�S�@��U�RF�|xo,�/���j��[���5r�����?.��^��|̃���|�ҷ��ߛ�*cF� r܅EK&/ġ�I���-m��d,,�{��W.dG��4�5�d��5���z�I�:k��` ��^�=P��Mv�,�:���#�+���ن�� �Z�����p���S�t�ۡ��6�5�¶.�F}���>iu��	bj%.�u���	�z���r_�"d��n$:�^� �P�x˝�G#���Ev=�lF#R��CD0@N�9��uP�Lp�V�Jp0C5�����I���c��3S�rb�8k�0���ݞd��0q�OA���\Q^Z��[B��KLث/Ӣ5���1R�s%����^|z��aZ������ټ_���^o���Wa��͘�lFm�x�^8��b�Vf�.�������c|�O��M<��WN5��R�3�-�;M�ß��[p��U &c�0nE�zʚ��$�L>��AX|�+\#�����[VJ���6Z4IX���y2
�l�47�F�y���N2k{��"��EF�Lr��I+�.uXvƖ�R�7�8���-�L��1��m鴘Q��q���*4��1��&�_hFw�pC$)��!���A?ӣ�թwjG��m�{�� ��>'F�m�~��=��v���6�QF�M���7��95��T����+�����ن`X���{$M���fN0�#�	�������2E�rȰ�-*���o�T��s(H�K�f�G�t�h���*�L�(�o�MwH�waӠ������\�Z� �se�g��!h1D���ū�`x��w�1{{��_z<S�#��=X)݌�Z3�W�F��f��Km�{w��V���dSW�%4�˗��m\0_^��Ŗ�7�"*�J�^���(�;�e;b\�l�8�����D��3V%�1%?��)��1��)��3�dF$��Ϭ�4&T�~��s\�IpC�U�"#����o�M�5`*���?���{�>^?�Ňj��S�˭7���(B4����Q��z5qZ)�{���QFˤ��8������{A4H�hC���R�	S|8���B�'��mJ��W���<��a��[�d_��M�h!��=��>��3��*ZigY����D��ˀ_P8[z�kŻc�FX�ˢGum�R����v�)�����R���m��P��R�q����96N)�0Jά�<!��)v&LQ�G�`2.�o�����NVuƞ���G�u�
�`�=�_����F������:�5O� ym=7��Z�]���K��n��Hv�c�$'1c��/[���#�f'���V�l�������3����P����Kt6l?��p����v����UC�l`T�8ʫ�D�ʲ�1s�nW����/��r	 _��7�{�?G���کJp\a��0*tHC�i��s{
�.9�BQ0ּH�6Q�䑯�i�u��3R���b�}5H��l�{ۇ4�3�����`�.�w�`'o�����sn���&��й���wW_�ϗ����ʝ
���W�#��Da -E���8 H��H,B����%1�C����\�N�+��j3 ���z 9�P����Q��mG��d��A�Cc��9����ݮ�� z���Ed�J�II(�J��5-
"퉆щ�%�Z�R7M`%��fPU7O���)�y�$�U�j�������@�F�t����k������㧊�C�QRH�,P(�f<�b���TL�x�U��Ƿa=�C|=�O*<��-haX!g	����V�6�m#>Q�p�G�� �T�;���62	�(�����f��Y����-��������^���dU��V���R�)�'W��]jtZyX%��~UL���J�0[�&��9#��J�R#���*��w�d먺�&�
�M�o�����ċË�ߊ��l���։��& , ��$�R���x66.�wZ9���*�7Y��$�ٳu�/,�F9���c[�K\��g�u9u!���!�z>���1SI���l�����*	�im��M�QL�={�^�4Y{)sU�2$��$?��[�gL�V�FJ��~2��ܚ�5��'�4f�s�>�b4ϻi<+��4����v�|��`������\����ڻ,������G����g��u�����yt�"���fz��vZ�r�N��<��{��gқ��l��MU�L���$=^���e����U�|��d����ݷ%`w��H�L��*�8j����'����O<�ݾ������ ��$�f�v�Q(k�z�4�
(Ot��Gv��ͺ�)�3�Y3&UY7�8���ق��6��RK|�~�|'+bd��:3��r�I�>�y!�w~�|!�qS����2M��g��n�$/�7�:�B��[���V2���p4]�Ɂ�\�����'7=T�=�W��A�D)�"�?)�U��ƾ�}����Ӹ;m��4��k��!��i�L�[7�C��K��@�� �����X�^$׶3���U��'E�����k ��3�V�:O�	�P���Q�����K��������~���Q`&�A؏+#�Iiӆ�Ϯ`��Y��2l�D�2�}0��j��/]����<�Q��!�$�4��G�f?�BK�$}����Hs�n wP)�p�u]�Ia2q��>���1�kfmj�G�/9��)�s�"��=���Z��N�[���9�I]� �����(����;�楪�v'q�jFf3�#�oU�%�'�^.l�f�
 �<������p�6�'�����[z������ru��͖����݊���`d�Fxy9`��X����ևy7c��?q)m���!�9����8^�4����J�~�4�`����V:�9�_��_t�y�QbG}<����;���X�+N�z�`�g�=����m����a2�8���F�p$��̂�>7gx?�9�*�	�����.d�r���2sb���|Cs��Hyȱ���x�}*@�~V�i�GvM��t�`�>�W�� ޠ?=7E�B1�pe����2󯌊<�s���zhL�z���y��!�j
s����f�d�D?=��̚*��:ۿ=�'/��z������ș	
�A��ﳁZ��_B�_s���(��+���R�K�덴��m�6�㪇�4��NQ�^f�b�[PX#�H���.�M�N��P�F������Oѡ�ɫv9� ۺ3eci��_�*0���%U�V��:�4dVٓ��a@k��a���<$t|�����Z�����k�C<���[ p��3�����VG���Z��i�.�U�O֗= L�N����F6��G� �ˮ��a�ы���w�6@����Q(��%@�yT�qFH/$��("R�X�R�M`���<pFGN�k� F�v�����<;���Ĳa ё�7�d��������R��h�L�}۲9�]��[=��lX�3 �:�6�u�U��Kn���_��ªq��h�
��"��/�:V��O}�l��&��q\m�������v15�`)r�Ƀ%c�����oJI� <��?)���b��Z&���I�\M���ɏk�n����V��e�5p�Z�h�V�{�҄��U�f��=-���8�
mX�)`��X��uy���'���n$g�4�m����=z�lc�@F4��s�V���=��(���t���S䤟��c��Q֣o]�aP�X�:Z�������اn�%8"�as0��y5n�r�;�q��k%Dj�,tI�֮� ���zkT'���o��Q�_����S�]�$7ӇYM`V׸*�q�'�:"���N6.�7�׏
��eŜ�AT����U�Ƕ�����A1lYGN��Xܖ�T�c)a��q�V` ��)?R�^�a0
)� \��)T	�E��Y����������UY���S�"t$��pNmԂh����/�T7���k^�k*4i�1U�. �$���L-	;���d+"��GZ��.�d#ƨ�/Zkj=�&��J"��.~e�F�? ʽ�I��%�`J.�c���Qk��[�݋͠g��N+[ﵞ��W���Á8=�8h�X�0z�3Uk*�{~ꪬ�R�rZb�������Չ�v�Ha1K��wG-����g�Em��z�a�4�KV��q�B/�
�Bhf����$��+)�v��8[�lJR�%d��Ju$�9��q� ���n�VY^�הaǵ�?�Ȱ1)�n����b5�z����N���.��˞���h{c�Qhc_���x\"�	A�!.Wܚ=f��j��<߹����O*��֘�揨P�ߦVC�NK�n@ [�dm7-�T,c�&��MY({_i��( [�*��'���E̦_��ʌ��/(P�G��a3q�w���)%Oֹ����)��P̓$Tig�e�I�WX��(�L��d�Dج�k���xl��L����LkVԬzN'����ޛeT���V�`��oR����e���v�4r-�g�χ���V�� *^d*pf�YD�?��G�+hzm^�*����rѠ�lI�̅c���i�Kv!U���Zd�4�_ �T!n2n�Fm:x�2�A"Vi"��̑��aL�@u�|��-h1�s��N�X-�f� C����Զ[�V϶���,r�W�&br޿�o��>a��p� �-}�s�D$Ӂ>�k�;�����ꑅ��%e�K�_	�y����'L�B�Um,"��{@{m��XN��Jv��HM���xlk��,Ά����<���P��B`�*����נ?�f�w"��{#��y�~�U��,Lj�aB��K�� ��B.P:vv���p�ja�HKBы��z��mo��R�i�$o7�hei=���8%�T΁
�y|Z���y�~�V���R���'l�	�V���r�>6���t�zr�����ի�/B��J�	���N�Q�3��5�ԯ�R�Lb-Ι�[�b����	BU<d����r`�)�nA���Ǡe�Kq�3���U�ax�;9gK�!Œ��'�s�3T�48Ⓥ ���߂�]� �@J����+�霙�#=t;�2;����Zw�8l� T���~�:̂�YuN^����H���|�;>�0��N5��<�̏���X��tӫ�k�8'�`���)-2�'����RNTG�t��j��r�!e5�rG�\��ge�uێ��AG��#Ngf����o,q��F���я�k�_CE�,%³h�r���&��Y��|�5�&��pQ���/JC�/؄�@�*j�^4([W��C���O�гmSz�ha;@s�fѺDN� (9���w�0*��R<�3>9�j��(}��3C���2�l�*n�<�e�$�Oe�f��Ag���4�qHA�P��S�����w���OǗQɦM������o�裁�B�[�FS�>t*�͡�����Z\W32,&H6���y��b ?	}	Q���<��rg���@X@���Ԗjs�,���S���Q�O����E#`���̩klz�� �Z#	���#s�s��r�o~�hH���O0PB�x�
c�Q�֌���)Ne�M�3�S�l^]ф3(��HF��NG���OW��� �j|h�z{׈D$�iz�8���1�f���T�?Ǻ�M}i6�Q����)d��Mxdv�D�:�*j�Y��;W��BPƓ���з��-��vd�Y��S�L!�x�5�'�ݣ�	A@�� 9�F!C�yl����~�=���K(�0����M8
�k"{~TB^қG�����n!f5��o�\�� ���F_�d��`ߪ�C��d՜e7~��ή
Ȩ�j6�]����-ؔ�+��f�۫�I�3��tW�@�&A7"r7:.����)N%U��v�E�׊�����&�W1��S5r�o��qI��*��9�5:���{�J ���d��Fq[q�+څ��4aeRt	���:�_�>��#��������r�4� ���j�?��{�� (�����o��/ODâ���,\"0a3�O\�����c|� o�Z}�M�.?n�E �)���JAº����ͺ��{�Tw���F?��q4RA@�Ņ�g��1ujq��CKYSۢ�G��Ӯ�?E{�1�:���E�>{�kN��� g~9��lQ�����~��%��=�ei�R;�uaf��O���4֎h�8c�gA�����0	6��V����6��=��WմS����������k��v|E���4�x�O^9V��7 e�*�{���(�d�Â�Ʊ쬝���B������d�W�,��i���?�����r��r��$���(ۣ]��oܭ�ar��',���$�(?��g�ک��^��<���sV���n
UUh�~����7ҥ�wcJh
Ee���W���u��	g_d�	'B��z���]�q���3�u3,ZJ�[�2'^a�����M,CДs, u?ˎ��љ�������ęy��>�f��Fm�HE}Y��(l��/��PҀ1�#� � ��"�tr?��^]���-t��@1v��mEU�ujr'�1[�rZ�95��w+������X�� @�@w�8)�p.�\	p\�T,�W��S����:����/��(���R\RPر�7�6�y��K���A<rE��fU@�Gv��jቭ�>�̥�j�}��T��]�E��b_Y����;A X��0��7�3k�G%���1ֳ��G����s�gvx=n��l���d�/�	 ��x�i7A����L�3����}
34&B����?�o�����r:c���i刯��C��o��Ĭ:?���MyL��8@"�*�iW���ﻁ�	w4���I�S>���F��u]��i���5T<<�H6���C�4��Vzs޻��9p83ύ�k��=��*�*����]^c>�\���j����t/�S���W�A�n����ޚ�qp(��}_�P;�ۀ��(�aHĶ�]��&j��̋o���q�Ԑ:�g��k�E	tf袪��	0��:�1�D+��d I�qO�fi��n��V.�_ҍ��DЅFTub<��W�պ��닁\�Р�f'�y�O*�F,�%��1��u�'�/��������,�f.�o*�:nr�ZB��\�̯��y:��з��̛id�c������}"�v�Hš^\���2��ADU=�c��$�)�*��H�f�Y���Q�0�_�r�S���Q8�=%���KҒ�";ޙL�B��
��zS��!��u7k C�K�s�逸]��L��i������R �����)��Ъ��c8V�9�A�A8����3��<��r(cT���$�:������� ���Ag��ݰ@��V��O�)�X'����E��}�Ҧ�9@�
e�M�j�n!�����y�䆅��9����Ae�y&+��coP�9#��f���S���NĹ0�ju s
q�j\舖�7��U���E�՝<�_� �d�T�=t�{�Nc��I8b{�>z�VI�?���߃�	ߎ`"�Xe���.:���6<L�F@Tmo�S3�-8�{ǋ��ė�^��v��+=�l����M�A�@H!�&S��$) F������c����X��H��К�ɕ��;s����b���:zT�CB�*06C��eF<L�,������J�nYƹ�yW�3����o 9c�=~b��W�)�e:jsE�=�����]ɗqS���"�Mpk;���^�i��������ҴƾA˺�7j�b@���<�)����t7����o�g�c��^S��t��q�Kh|Fy�!#�����\��BO�r���7b�_�^�#u�K$�coX3|�9�W`ʖ�gt�P7^1��p������y���:窆.�6'$���3�����uJ���Z�c�����됯��6�H�t,g#�.\���1��k�r�7ʎ��VX��W8r`��	�!��Vu���*�!袪��l��ygf܊渧���s��m]��8����lMX����J�;�0Dx��y_��Z.6�U���}n���ȼ-�ڃ�%��C��zW	����(�d�
!EdI(f���wz����؅!�z��X|:`CK6��{���t�����g��^��*Z�������FU�\4Ѧ�����������Ք��I����F�ĩ�dVAdύ�B��o�dD��'Ҏ3��q��%��>o�ϲ�P�]|��9���X0bY��0-�9�TM�����y�5�9@]�Y��&~�F:��+��#*@��?�oh	��#)�r�k��3��VZ�s¶ɶǵޱ��+�z�.!(u��E�;ZJ8�-�=+ա�NW�$�s�@}H�!ݬK��a.��N�7+Ł�d�H���#��ҧI9���l�a�3!�}-��yE �L'���&u���p�T�a����*	��8+����:ύ�-`r cH��ڷ��s�#�e�z�l�AtyD�K]�{�����ё���^?�y˺+"܇~H�F��^w��3�+�Z�x.c���-�uR���L� �qL���q@���� 2X�������ZbE:u�d���2�x��~�D��Ri��p5b��hV�~����J�*�V8{�lߵ34R��D��O/� )�l�*�����s3!gZ�(M�P����Ēs�������}_V��N	�Rc�XN6ڨ���%O�.�-S����-���/�"�o��W���
�0P�2�Ü�cˡ�����|w>�]2�K�D��j�V�9�2�п) �p\nm�~%_�(h�/l��q��e���a%N:�5OK�Q{����Y��%ќ���Ԥ�K��3/�B��`D�������S�ӠX�vy9����D5��шO��V�A����.�����?)�t���?R�K��V��I22T�N[%mY�@���>��D����Ңv�ի����x�_ְ�����t�;�Tդ	"L��*/�)@rr�^ٚ�3����NN���kc)�f(K�(~�7.�NW�stc��B�=Y��\��	��~«V`g���k�}*R�mPj�sbή�����5�k^ �$�,�U3��%�i�u  {"��c&��w�ꝹJy]��<J�0���#���������M r�5ln	�~s͹�IW=%[TqRJY���;�ϗH�R�le�$��\x�{I�Z��cdE+?fpQ��%���E�Uy�+S�_)C��)�TF=�"�&5���:C�+vx�̂)�Pg9}�Kwʺ!|�p�q���ZCúq�3nXD9ɸg�۹�Y����u(����qY��S񻠞H#X6^C�s�g!��L�o$��/�R��e˷�]��n��a�J�q��Gk��h<���j�񊑺5�1#�E	�֦���Y��a����h\2�����W���vJ��w��c�DC1��<!�Qgt����*�-�|	e!A����պЁ��<;�#��Z�ЍQj,:ԺH02��Ў^�Ƹ�.�|}S���6m�C{?���F&������[�i��TG(�M��t��t�xo�h,_���{� v��5�� #<�3��5_C��2��� �����o� �������%��e������~ү��c�lK��5���9(>�0�K(�r�g(W��<�.=�P7"������4Ҧ���5vC��F 4��]�R�9s�����}�p+y����J�X�}�^�/���k���6�0@iH�|�ȕ�� ������{^T	�֚�1klAV���Cmx1ߊ�T|�R�.��~`KIVM��G�,f��l~I$�>�T
��ق5j���CC�*:d��6O\�qjs�!�|-D]��\C�D����"5�ʊ*R��oX��I�g�G�������W�p���1��bP	 PP�����a *Du���� 3[�n��f?sO��Gȉ�M۶=�N��ƕ8�K�b��C�^n�
J����H#�"��͚��(Y��%_��qSQ�T��g]��]��Q;O�3�Y|���������FaʄHL���
 �h�)f~L���A���u�ǮY߄�E��!�	CH�
r����v��A_�s�O@���r%�5���ߘ���Ƞ�<$s�f�(���N�T�����O�!�
9�S�^���N��Cw��� oe\3�x�!�U(�')^Dؽ�D�^=��h����8�w�+!^@9!��?�������xڿ�z��!��c�K��+��!3�z٩s�6�!^��H~�r�v�Z��~Z�u��)=��r\�v6@����WK�����gs�_Q�`ˀP�2�*}�Ս!A�L�waN��qD2�7�m���N㰿[�o̳W氮�
Z�_%)߈��k�v��l]
��FF�S]k\&/".���ƙ�^(�s��4��*ű�/��Z+�y]ߖ�FƐue!�ql�#��C�մ�� �����!�?Ԇ&�a�W�����~o��r�l� ���!�U�k��b1K]A0��`M��K�=�0�=�6X�/(_��1c������'���[7��C�������u�R�#
߂>�6��TkZv�ah.��m���|��*	�wA� �h�tX\��ۇO�Ű.���R�.?�S$)G���[�:�B��,���ƾ��
�?<��D�ާ�-r]!c�����UI`�y���>䢖���K���w8[������P��i�΃Zy�W�4F�`��k;3ƕ"`��u�S΅��u�v��X��wZ�aKSUL����v���*au�gk�/�����3���l}��cl�X�K-�Ј�f�ell�Řvh����K� }G�7���(+j�c���.�����hT�4� K��pI!�,�y@|>��wT+h|˿����vp*o����A���aG��JL���iY�9�[��p����^OV��ߜ�I�6�M�p%Ф6�<m�����^X �m���Im�EC�3����DƶS쿣�̍Y��8�#` bV!��7��I�Ch�l��F]��se{����n'V� ����e� ���(S4�����ۊ=Y����o�3?��A~G�	��7ߺS���R���#E����a��_�A��{:�NDH~��|�Ϧ�Ĳ���n�%^
=ۃJ�� 6��?b!(��j�h8{�(.���j�u����p��٘����"�9ݷ
��:�~q��bӞ;q"�w�-���bi���M�)��\01�A��@R]��m�2/,�Q�tS��)�	7\�<�u-A�p�D���ۗR�ۓK�lv�wa1yT��|?9`��:�����ԡ���EG�_r(F#�`�9(�ǒ�����X������d��������6�� �[�/�n�/�^Bw���J���
y�����s7�Q�U|��e�1f��S��B?�h�B������L��T?�g�i¹ B:/d��\�Zb2�@���fe`���Sl�l�����O�~7>O��X ���q=[O��	�G�k���V����_�߄�2+
���6}јճ*8:X��wrײ���#'��~[�Y�u��1�t��.��;��{xe�Ȱ�2�6\gR��$�L��n[�QH
��G��T�b�'��.��s�rh[i�H�V�����i�m2��
�H���G|�K��v�JH�������
�J�@���,\�H>�=�?Dp����o4�0�
|j֖�?�:���|��VOp%7�In����]�Z;ɮ�Z\h���h���l����tш\�=�hb��sU&��<g�s��P�C��,�X_p����$!y,QO��'"�		�;'�޹�C��x�\;o��=4���U�h����È�)ԍY�>`rt�4�Gf-��<�KW�n04mi��2��l0����ԪI ��K�R�j���[-��9#��CXx��ig�dx�>O'�GjDk��@B��D�؉��?�s��(��M��鮢�ç�|��2�{���t��C������~�����l�E��2C�j,q�8�  ��2ԏ�5�X��^˸�Js���f��y��[ř�e֧I��eX��ւ���!�eM]eK�:�#*D2�*�	Η�6PR-������c��cŀ>Y�<�5�v����u�V��'C�RZ��8��WYݾM�3u'�����^��5su�?�ƙE��B����\_��L�J�0�+FA����0ՙ���|ҵ�_��Pw�����WWj�7f�kM������E�䄬�"���2�W��mN�U�#.���+o�²Bԩ¡TX�BwK�ж�v��7�߷� wR1�p~��
�j��������H��K�I|������ƫ� i���31�e�u��GL2ңG��qᕢ�^�$͐k%}R��I�����V&�Z
뷛:�i3CޥD���o�;�*ov"�K吒��W��-U<�f�r�8=D��]`���5!VY.7�A=�ٟ��!PZ��^�?^2��$k��VnH��?y�
���	���Nx6CC�V���\�>�]͗�x���Y*k�<�|��{~�'e�o��8��UC�䬋�jg���I���<V��'���\T�k!s.?+�?)j=�ͼV�E���V$�;i�mryk�қU��U�V
ٷ�NY�h����0|�e�^/��	?$#'����h�_�.h��A�@/A�!Yײ�F�&�`��9�����L�#��S��ҩ��Y1ʾ$Y~����O��uS7moO�1���a1�E"C��BDK��8��u^���<l�)�6�`��ot�� q^�Q���5Xd�7��T� �S��ʗ%��6��)tp��r5�F�����wx�����1��6�����j���!�"��d�0k#��v�����@�9@��zpPfV/MYNt/��!��y>���zk�������p�#�]��!�R���SkO�N?ϥ��H��΍�C���� ����JMI���g�q֔�ߟu��7�F[�|�]v%.R�%v��[v>I�!Z���O@K��t��:̍�n�����7Gyw1���ͥk�
�{�vQѯtQmm*_ύ�)r�"��]-��Q��W}�U
L��Li�t ��
��[��t^sr5�Б�eq�j �W�詓�W+�]�(_R� ����X��]B���h��r�ʉi��:8�)�:�qm|�		~3�Ф	��dÎZ3=����� �~r����=�j��A���^��h}?�}M@�ܣ^�l/7ʿP�튞��O%��܍�5�b����$F���%�_AP�侷����5�n��M%��=����?��UcY2�)x�0܉$+�$؜�fﬁ���>b��C�f�vF�$́	����@�����P��#v�LK��bJ.�V��>�j�^��Ъ�œ]ʤ-���*Y]�-�w�[H�n&�R\+ ̛�?���No�(L>�0`������m '\iEg)�"�~�Sp��D��_%n����W�(;H�h1'�;�𤋮���>��S��˚��L�ĺw�+��]�u׌aNG��o8���>g�Ɯ���&�mY5���i#��%��
<aMU�xS�ʉ�$��-�m7A[y�H؝R��J����ɡO�o{*����V�N	����
˙HĂp|#1ȓ�#�>�pYj�Qr45���_�Ƌ[O����8��7C�:��)����9^bj�>��,3D�3�Ͱ�)��&\�<Dc��B�	��F���nt�@��,�pY�-"_ŜV��U��@�֧�W��;GpR��JF�4�sU��g��-�����9*�;JڿQ��~�Mm���g���<.��.��Z��x+9��@���kuŮ��8Qu���˙��@�Ft��<�t��bv����у����8Ҭ�,��QM온�Ʀ�=4��=/t�k��`�Eѝ�X�>�'�����ȅj
9�Z��(�1�|�<k'߫�v�5hD�9B�h10��ص��gp�L�j:
S�ƃ�Y����p�c8�Q�[��>�$�u,Xge7�T�/yֽd�\I��+��H�������-��������o��Z����y�TlO�����6���|D6����aC�
�X�w�0��
����^6k����R���,��I��c�U�ں£_)^\����-K�C9T���QF�E#���&��P���l��6^Ua����pgKw�T���Iz�VpY�Z������Y�!mU�S�~��� �͍Ur�iގ��>(}r�&�k��+��d	� ��=���b�ӷ����c���)@榿D��8�88������a#�z��	O�׏��WĞ��|���wĽ�]KI��R�'�����ߟ}?��,�)��x��WhQ��e-��{Rl�#Q(�P����J�e���X�&D��7��g��Р���?��Q��K����*�w�,H1��J>d��֚R�bi0�~���Ւ���Fn��'�-��~���լ{-�_m��vE�i=�T�:x�1��T|��+ǅ��,>Ts����\)���F�����6M+�M�i�;�����ښ6T��.wPϕ�*4p�&ު뜃�L��2{�����=���S��w����i�ݮ�3UcC��!H���f��-x��2�3)];[-����ne:�=U��_�X؃��肯(�6�/����B�]��A+'M%q��A�g+���q���9����[9OY���`���
N�W�凇��Íqڝ���ʺn_�?-��_ڳ�;uFUH~� ̷떑o�a�r�2������� x`��=E���c-q�r/�X���y[&�#M�C]�w�qx\�0W�K4CW�����Ɗ@)E�����Z��P=��-Kt 沖��4f��<}a��������HDr�n(�5�jK����Z�@)O�40b��O eOP.�1��Y�58"�%�ۺ��if�ή��ЈJ���V]�u���(����`�lx$�_�}�&�7�[�W�<h;�����!�(�Ѥ ������N;���D�o�C��
�!�<��8�&B4Qm	��Z����1�V���1���rѷs�A�B���1$4������J�XRi�O'��JB֌��7�]�A�1x�1_m˽������o��u^A�p��}�5���P�e���d�o�{<(�V 5�0_u�&�H�/)�4�A����M����ƙ��iNx�ʠ$���0�5JP38�#k�:�_論�aI~�mfDJ<RŃ����ɓl�R����UK���K�5�b��F'���b2�fT�k�3��H�}���}K_4a{�w$a� �2a��S�[��.��T�#��k�a%���S��M���dQ'U��|f}���L���ECX�x���<RȲ�^:����o_����7���1$��  ��w~=�ޞ*a����Χy�U/tm8)�d"�R�-ǥ=���a�h��qK������#M��j`�Of�ᅼI��Tj��Ľ�r��Ѓ�1�l6	��W��v;@R\s7A]׸+��좕�*d0�'+���ƶ���'�v�Y�.2�5����|�\?w��(�Ł��&�e���U�h���T@6ShL�4�E��k֊�~��ws��5��GE\b=� �ŗ�7v`s;{�M&a�6�T��l���T�j�dl+;�l`��A����,K�<\���#V,����b�*��b0S=��2���������A,~#���i�x�8��N5�� ���%��5�	�)&7l���Q�C����Q+����识I
��`�����4+.G��b�w��+�D
F,�R���G��+�:���Tc��_N�C�I�̤�� A�̞Y� ������䲊��:����3[�R�'��}��Q�P�-��W4�E8J��*GC�yV�6�S��z 0s�=�;�� �����T"��U[U�Y��b�"�iOo�4���T�N39`���Z�J-@��x��Y\U�C�������5��-�����=RD �8�{�����ÙJ��n0�ϫ�U�m@<%蘞�	�Y�O������Pu�C
Z
�"�?C��b8CVH�ok;'k=~U,�1��V��"�S��6K����Ǉ��.-#���=���[o� \z�S�/�J�"�*9�}�'�<VW<7�����ݜ�4f]=�����}/�#y����hY���'��ҕ�K��k ,Ξ\���M�c�,8��O�j�|��h��cL����R��s�r���	�5���̔1�q������0T⇶i�?W{�~C�$��[��m�+��;)n<L�1��M�+���ȃ�h_�v�^@߮%[�v[4u,���e���+"���/g�M3ԸdYX���?
���Y��q�Y%�,�R�Z����	A�i���:i|A���bP�A^{�9��+�V��0�)_C��R��[�zL����ܕu�>Ah0�����M�2���=%�vt�.���O�X��WŻ[�V�@�D�7�?�+�P�У�:��T������I���-���`�_M��G������`�@De ���y�M�{�5~eɖH��'�Q�I�]U��h��HzKwc��9|��@��bfMzt�갮����v�RD�2?�����ڗH��<]�J��������|�oޔAz,=����=�ݽ�;0/n��(ˣ �B����=��5[�pz�l�\pX�X���II���sš�y<��g��6, N�����)�
�yk�ݩ�r�4���?5m���G#�<�����?fc�N/g<Y�EW3�t�#�Xz����V��z��?��/y�PІ��
-V8�o�S��� ��� Ùy�o<е�.��Яw�$ȌW�5H��q�}��"<=�������_7��e��dկ��1ߍ�j�;�o���{B�Jb�Ҏ����;h;��:��L@�b`Ƭt���X��@�|��a!_���yղ�AfԬ��.I����Rwރ�o�t
���$���.V�J�^�� M���&���b�a?8�ɠ���$��D9�$���!���UB�A�����4[�7%(�����Q�I��	x۝��J�dAy�3Y�������es���b��&���`l����YC��o�OƯꠏ�{U�%�E>Z�!�v0�P��Ie��⫉DMr�k�e������t�q*��o���!	k��R;�c��͇}Fᮼ�IRm���ŗ�0lIL��)�V�L،��E���X��;���DaTH�-��4� r��=��$ͯ�B���i?�A�[/��S��Gz��u���B����;l]��ʉ�fT�#c���(�@���T���3J@p�8�[o9w���v�H��C��3ZR_Ǥi$e#���k�H�2���VN�0�� ����Τ'�d>��3���Q5ťG^��~1�y�O$2(����{�����w����6��I2��VUv���p��M�M�� �OecS�ec?���� �%�q1��ǫ�9�IE� -�9���'~��6���:G��'f4�������6|`Cj���ض+"
=��ݠ���dݩ=��đj2V�P!!�&�<���H�s��&��&@|�S�Z�Z��* ����viC�SW�q#N����_#���������R�u�ᶚ���+P��w��H��ݩx�%�i|�ҕY+f�㠻]}̃�ۮ{�mr�=�ZH��(YS����c��êyuR_���i8#��-D�(N�aѢ4^_��7u�b���ӖTI>�볕c�<ԎH#Xf�+(��>����(>3�۱_��1I	���x�`��+�;^R�D̄�&���6� ��s��]�̡�W��?����m6}������}�#?��:���F�et�Hd4���7o�p�C5��"�Jꘀ��9���:� �C�؄��xQ�ү9<H'���DX_�)��@����L�ݖ��SG��c�C��%h�]���Ԗ�#/�h�d%�+���
K49��?f�y�5"~���5�(��~ͻUM����h��R����-Z\��u ��V k�/Y��]�l#b����q�-b�{��#@9������h0�N�~EOJ��ı��"�Y3��A�"���qSԿ�����WSf�~�?���BAg��Ŵ2p��F���ѥ��^o?=.��>�;U?�����^�9Zmc@:1 )ǆ�B!��a{?W�|.�*P�7�{����5-#�E��<*���Sl��i
|@��� ��L=�,�$�_>J�n�F�֩9���ME��hEJ���*�aI���"��\.͢��w�4��K���8��c�t�M�z��rY�k&f`�
o������-^����XI�N����&",�aV8�)�������K՛���Ui��ue��g_�*�w�pO�fʚ�{�:�0�Y�h>���C@zr�W	�BI��O`����ڙ�<����׃�:���r�*�;��+tf��j�1���yg�'x�$#[���V��rI1�	(D�B���R��@ٗ��![4u"Z�`y%ZXa2��K<F<9�8��=�-��9`2���g�-�h|>Y�w�Cc(ۛ\�r�g�}�2̯�rk���󵊆��\a�!��̻1hK!<���p�'qd��6��@�y�k�zٯ�;`���芥��^��b�u��z���sP�E�D�t6��l��v�(�_��U��v9yE��=��9���'7PK�F�%q�R����S*D�X_�L1t���]sLs9���88>�5^�@��
+��g��_�x��Y�������0�B����k��:>ۡ���d���� �ƹ�6Dy���v��I���ɇu�wt{����`�	�mM��g9i���t�p_����'%��	c���e	Ğ��߆`ir��w��\��^�T�XK�?���`k
����o΄��Y�7�$���h�!9�Y���[[;��WT��: -,��Y����^*�t���z�IWX TF鬏7`���y���kJ�vL��� �4x���,|�"����=f�
ʀk¶����*c���1��΄���+5��u�0�+�� �"&��3�Z��e_�D��E�zk�&�lz�˔^������(�c�^XF�@t�`���$0I�k�xM��I�������
��(�w]��K�B����6�z\*�GW_�t��bM�Rd����f䛠ҔN�x�`�R�]�g���me�7���G�c�/��ݻ�_�%E��׶4.B��/Ҳ}�ü�WJ�7��{��bּm~`�ƴ�+���1٥N�v�'���1�8YR����0���O�����tZ�G���N�Ye2���*i����tv��Ig8m|�U�T�c?y��p���D�:���į��?Oj��XI~v^g�)ފH��$2*��M`�y�Κ�yU�"z� <RY��S�A�X�j��a	*��Vۇʽ�2g�o�>�R���$ӾO$����Ҋ�p�Z^�-�F�j�L�a
���Q�G�ijz�˥��������o�r��q�C=���>$п���,\�	�m���G&Q�bӈNt{`G���y{�Ż�]~3u��"_�Tt5�T,/�=���ۖJ)Y8��t���Ȇ�Qj!Չ�Ѐ�Fд5��SY&�Ö�@�޹��o��I�t]o�0"E��+��|�Ė�Szw�ô�g��GI
>��d���F,��#Ẑ�#��!�{\#Z��ؗ&�p�{BQ��S+�7�)+]p�"4T������-���,�ֶ:�|v�Ӡ�E�|?G%�yR�+K�S�X�֝:����܁9H��HN!���Fw �G�/�L�>�޲S(WL�����s����-�W8miVo���olF���@�X� gV)�J�2����$�~3
�hY�s��P�˒�xb����c��(�o}�;U�S<�0�(�}3�:F�ć:c�3��'S-X��a�Ti
#�`� ��L7k7~,Sb�E�jE@�a�C��q�����D�T����)_e�1�&��EMDi0���V�%w4 �u�Ę�2�S�|+""D�@{ewz-�c��Lkk��	�fW�N]S�0�HHÞ��H^-���S\���[���4(!���� �U����De�^ �<e��=SC��~��	�>�A ��MH}K+��T�/l�B/ڑ��J��"�91�r�2������$MI�Ӣ�Z^߀k�e~V�6~�p���yl�IC��T"���^�񷱜�,\	M3,�V<x��%��n��p�Ҫ�\sEM�Cӧ�G�2O��+��\	��$O�d�E��+�J�F}���3�!��	؀�nHUᄾ�Q���W�|;]'k,an�W �K�hU�2�aI�f����J��n���Σ��3��fo��8S���2��e�!�n�е*<���B�-�@���F]0)����ۉw�WX���ޅ�{ϸ�B������5g��Ck߅�)�
�pn���B�a|�k��6��׈�du�R}F��}v�T��4H�x0N�y<�'��>^W�/��˼����4k��(��#��������7��9�k B|D�-������*ыs
C���z�T�Bi�b1�p"T�G8�lэ` ��������V-�y;l�A��9���ꪠ��j|�۩¡�E����,e��4����ac�ꚃzx��#Xj��~�C	�]��b��YbL�_����{�F�"��t�%�-���Y���DA��8��>�Ϥ�݊J��G���3���Ee�8�0;*� ���b���_GN��<�ŃL6V1�n�4�
H�(�;X��Z[����q$�k���U��s.W����N����4�������Gr*��^kT���O'�X�Le"R�i 2�����>��=��.�o��� ?+��ݻ�1���	:T8i�4���a��2'�{�u�g0�;ޯ��L0��_Y9�Ƒ��������O��%j9sG5�Ϧ�WE�Y%U����ܩT"	����]�:ۦ��������_��jaD�Z2<��+
��nr X&-RUk3g>}�v2+<IIV��l�a;}Ij�>��F�W��^���L����� ŉp�+p�oaJ/V�U{i���m|+j�^��}� ��^MT�=JQ��!�N�~ȱ����s^��B.������u��l�I��Q�������5UelO�"�諿���Wm�5ou��_��}bq��_)	���<�pɒ�W�Ƅ0
k6��7B�`�X�K��X� ���QV1���Dr1��F���Y��u�q7�&f��#'�M�Q�p��(�+�����Q��4r���m0 4�2T���S�x.χ�2�a�R�+%Z�8;TbQ�E��l�����٫Н��M r�<L@�4R��z�BW��������I��x���\���D�2Q˻�K�h�ŒNf=��殊7��=|�%���WM�v#��uU~�@�9�3��C���
��qj�$38��	f�	��i���?�q�\��2��S�[l����n��ze�.|�T��r��HT�;h|T@�%�A4�S6f.�#�z�)	�H�ڟ�֖v��@ȍ��L8~!�g6����Z_�x���eT�q� �ď��/j2�Ј��)y`u�~`	��>إ*ٝ@�u\��	�@���N���Ed򖩶bO�5�n�V` ����΃�_�Q�[�'v9e�Ӏ){+Z���6uj�'Pr��1Y�椫��0Cۛ�E� G�Ó��X���iP`0��>�v�8�ێ^���$*��(��Xy���)�I� 	��âx5ޙZB��c04M��Is��51݉��=_]�#d�~)0�0�u��f��x���=��L�]�� >�b�8 ��Z\Z��w �.>�7���dwRZ�a��:&l��-��W������:�Z@k�(~��ЍN���6�w8�f�(�@8�.T {o��\;��M��|��s�y�M��!N��Ņ]a/���w�ҧ�E�)�����=�z��\��T@�O�7*֡��R9�2�-����f*\�.��oz�z
 �<W���f�V2�+$4�ц�,h{��BxNF��7W���r������淴�Ec�]*��bӔg�'�.�J���S(�J�HDM*��eT�%�20��**Be��KZ�b�kv%�߂���g��8<�<�hf�G>�c��%|�K:b�V��K���<���HM8ÔτƏM�Y��j�R
q,y�QDG��:-�(|Ʉ��5���<R:*���Հ�c-��p+�1/���F��K�F?m���1bYC �߫��^s(�$-Gܾ��`*��m%v��V��@�%��_h���������(_h�j YB,DM7���ت���+�C%Skb�â=s�:j��-�
�W�+��C�x�('<�	�|=%�������AC�z�y�[Feh���MP��u���p����*F�#�0).j��~��2'�����3��]ۏd>�4 ץ�M��A
e�ebU!9�x5p2��F�[F��Ƃ��(~�S�oJ0p����\�Px����q��;B�5o�4�����n�ŉ�<���ʝ�7���K����Nl��耮�B�W���_cK�M&2asdp�bsW����,Z����>����ls&�K���g
Eu���b�=�|/�����S�������*��6k���6P!w��碨�	�4u���l6�������,�:��V>j%Z�z2+\�tO-np~�,@X;����nN�c�{�Tq�
�=A�����rlE�����H�������>2��C]�'�u�ަ��z]��]��YؿV��pCU���(}��'֖�\S.!\i1�}.@ѽ+cr�*�BЦ@����DVP��jb����J�֋�P�|������PR�X���$}��B�%0�� +L��0ڼ�̧�-��7��00L�b�Z9�"�F��m���1�} �лl,?��'A
�dW1��d��Ӛ.�P6j�d�o�r�ք:��D,u��B8�暒!Rߵ�2&o��sg��T��[��p��a�5�#����A�!�������?̴��n*:^X�I��Lmk䚬����ځ���Q��T���j�8��� ��:�9�E�c�[V�K�$������������g����{a5@�4�_o,<��Ѻ�`4c�G�]ܾ.�����u�&o*�O�E���o�6{U��M��wU�ܸ7z��b8k��MN/󖥉�m���I�--�G�Ҳ��9�%�����B�u�h�v���ݏ�@�.�ӛ������~agp\V���Dfz�T�}�������F�o��j�u�$�������(��
g�2�
�MQGa-��y5lR�U;����(�� ��h^����C��g��Y���J(B.X7T��L!�@~�O�0�<�5�>"���!Q[.�,����7R �����KA���[5�����0�� � T-1'�m�`��v8B6����5�
0�E���;����>��
8�.Y�ǐ
8d�D��2�l��x��e���T&�9ވ��; ��#����#�O<��S�Q;%)�u��Ϡ	L7IU����,>�:	��8�)��T��ll/F�_�k���~ݟ���y/�4-�WucEH83��<:����zj�m��_[�:#�ڄH���A�0�E��#�������;�PW��7�v�+����#X�9�x]H�� ���g6����q^F(�l����磂
�Q/����å8H��GN$?��[�z�wۆMM����Ŵ�5��������%~[|�K8M`���}$~�F��G�_�K=����J���!�%�*R��6��k[��=J[��$5�I�7P\ۗqi� ��$c�k&F��k4<���Y��n�S���NC-�������I��G�a�����T�D(P�ʅ��v	P�
ý��R��>if����^ ����[7Q�v֍p�hUi�Y*�.	'()եҘ�S��P�z���I����]X�������Ę�m�*H����ڣ��죋�FPB�H��PS�/(|/x)`o�|C�/n�Δˁ� %���Le�8���>� g
��6r�1��F~�o���%^��
ʧ@���`�!ゞ�3��g!	m�>���lV��~�y�!��W���f���{�3�C���k�f`oV��
:^���5��?%/
]�t��!��.��l|N�П�m�0�ݫ���P���:�~�7�EoĿ��KY_Jl�:���{���%h��E����(�P�E�M�=��&- ؇ڪ�Wr�~���̓������������H��@ԉm�0��g��2M��^��FW���:��d�{�fE��p���Ǆ/%�Gu�-9��yu9V����0;[cs��x�d���U�@T �L�|�;SvQ�3̇P9�K@E��藚�u�u���X3_�m%��uB�x�B��[~sN6���x��Q�e��Щ���'K�A��Q�`GE��lq�$[�-��%U��"����ڿ2�>����O���:���p�|��s�6�ss�g=���Q�~���K�'�p���xf�"��<'a�N����Y,�b�j�$��d����/h����0ֺ C���X]gvL;��!o�P�DZi���9����`{�@�\km�p��~��x���bvC�����c�XF�?eP*���=Q��1�(�L���ۻ����V�b���V,��F-��r�(�L�\�~¡A1~�m������G�ʬ�O��r3N�7�X`4�s���)�
9��t�YT�9������ +t/���InN� ؃@���T�*I1���uSc?t���I�RԒ<~�n�>B��!X��!��m���c��a4(U.G[��|U\��?
��!�L#3i�� 9�&��2�@Ts.����?����b��exL���h�Ho����C/22�D$ �D�q��/�h/Q����&B���#�/�0J�Df2#S�S�n�[X߿�&��}8���9�'��F���^z�q8���f�W���=�1m�X�Ǥ�`�i�>�F���!���H�+&9`i�nAbG8�׈k݁;���>�a��������ʎ��j�ކL�P).)�g;�5��#bT����א�/d�V�|��U����p6�OԼ�����@>0:�ULJU��G����q�U�#��"���钋΢���T� �q�2�A�%�!P���tk��X���`l�3-�Z=JLS#uL��x%�S�!�>&?�F��^��?�r�?KZ��?�� >��u��b�+w��n vo2O���c
���|4�u3I��^(��GՎ�6�Z��#u�.G�������`DF|F�eM����n4�����"��ǭ	Ӳ�H��DRZV�LR��nn��o鍇�lb��$E��?�. �V1eDC��@ra"��2Wt����.��m�p���I�^�(b�hn�u(یI+��GZ��wȪ6�f���p�է���Wy%�����@&ҿ�\B�u���i�l$l(�4E�ꇦu�����)�%�D	ͧ��\�wd�s|��T@ʮ�s���(�;e/����<U}1z+'����pʓT���4����@��  I���˄eOTb^��-XZ���.q�Eo�1���J�܅��BX#�^>ޚ����N�O2�+��ڪ���G�  p�����'��fI2������U�go�[ +�s�]S��t�h�6�1R�ZJ�v�MA/�`�I�X6�%�j0U��D�c��E=YA�H�1� �V�&ْ���s[���&-��#
����x� /`'�v6�5�b��"D	��M��9�dk<z�U`$��:��z�"&�X$��T��_�@u�=:P#We!5$���Y�+�,���n���-إs~���1�*
F�Yb)�!**��80�� +w���5�gg{�	�mM���ݿ��>�}A�MC��]02!N�w��J�pW���G_����1p���"�5*�0ޕ����⼹Pqr��z$��0#�>(�Az��)d��3CS���nS����4n��5�@��_3�Vqq{,ג_�!���vM�F�;�ϗ��nW���U���s�$Q�MD��%�Yg�����r�{O���ަH��D.��Ը��g�L��4�W)C�Mz�h���
��3�Y�X�{>H-���\R�~�X�0�+fi1��z��U6�V+.?{�R>A�@%�?�Һ��2����������췣Q=�u���L{���s_��4�7�/UFN��+�C�<))
�n�-к���%jvh�0���l�����ݥ&�h{K�Box�+� -��/9��A��s�k��ߗ�a4FkQ+�b{�Pb���d��.��6�l�1�lA��P��)��.��h�Pf� =5�t�ߞ	�'������X�d�^緐\��Ң[�vGsQ��#t���H��%��c���pU 4��#t�
�x0�B{}D���˷jǨK��� �j,���c�%�l�� ��j����A�Y�0ͫv��e�Ew�D���$h<T�fĺ5()գ:GGy9��%�l�&z��f�D��(4aH��b��!���좉 �=� �,Q�Q1���? ֕xA?��p��7c�*�JҿȺe2�:��젭$�C�H�n8�y}2}�+9�m��Eh�����۽L6#�E�I9uSŏz�U�Q�k|�(���_���`Z�Z��{�$��2�'#�{2���������(-a2s������Uy��1���zk��Xͮ�|愯�f�MKdyV�\X�ڜd�ɒY�3c������1,'��u{k��4%�lX���*!�����v�ZA&@�6Ҁ.ޠT��Z� 	�A����|�T��D'�K{cH^+��i�rړr���K�H�ou���[r{=4�D�$�gM��%Ye�6ac��J�v��ɸ�G�ޣʛ����G"�(�@[|\�h�8����6��49qX	�V�X%�I�Y�k�����.�:h]VZ�h���X2T���)���Z-�|�ltXN�/�^��Lɾ�����_�O��PO�w���-̑y��r #���KЩ;
�A"dq��f�t¨�_h��V���}vV�'�ċU]�3�*9|펱�v���F.���,J��7#���dP~�^\�o;���4�Ț��vR$�F#C��'�����=0���&�e�?�V��~��˙��틴������
�Q|wK��c~�	�wLD4�ҲyU�`
j�����q�4�w���_A�[A �2�k'so���8��M�(͢��
�?��>�e{�a�:H�'�g�A�Q��Z?µ����zΩ,^_&��2�"[S��7�B�Lz-�8�0���zfmeRHF5�U��Խ0���J��7��K��j�qc����C�;rzN[CoRt����J5�YO^��^��y:6h�@t�7 \n8ųTK��ױ��`"��x@������M���>���)G8�n�H�>�O��t�2�\.�~��\"_�6_h��)[�^����5>X�[�`َ������� T<���m-*�c.g�Ү�#ʠf��1t�Sը�@8�[4Fx�{�]�iD�l����D�[49q��3��F���_^/~T�t�nt�rWi��V6��e�6�tv$ز�3Nvze�����g��.R�2���r�NZ&+�*�lp�p����H6#�����m�'2�5�J�Y)�o�A$��.ծNZ 83Z_X��N�<��|�Y�V�6��jn���j4]�$3r%8���Z��( �V�՘�	"
%9 p��+��Ög�Fqսq�i����*6U���˂�(B��ڤޔc�_�B�fD�}�d��e�pH	{�8oJn�2{&�f�*�,_Ų�W֮��eh������j�ef��zD��p�PB��;3Jĝ�-��q>����l� �"�хLL�n��`�nm4Q���s�zY�CYm��p���W�ʺ'��U[m�e�l��je%�xY$�5�*D�"Ѩ?�Ó��[��5N��b�';$�ߥL���[#`�Pu�t͌����#�KN0��
�&{��Dn�	E�7y�6W?m�Av~V�v�������?D��tq�?��U@-�MN/�/+��tÑu���'��?j����6o��� �S�.�D��8v��������Uèr�X���ܩ��D�&9�N)�y%yZ����=�w-kx>Yxs߯��շޯ8CI?�d������j���o��g�و��]���@�	Y�;�S�+I|M��'l�el8���f5�˱�*�cu>-����]��wL<���<�H!�i_8��ᑈ�b�����}5�: I �K�*�4��fg3�~2��K�4W�R�X�*�٨R��^y*pW`��qa��A|����.�3F[�l�(�0JN�Nر9�]j}�U��Y�w��\\Pݴd����^)}C�Dһ��u��[!]*!�T]�Z]}���M8>+| 6MsJW�!�:pB$���Gt��ĵ�k�5�e;�o�B���>1�e.�V�d.ϫ�ƎyWY�h�	Ǜ�����[i��#T����Z\v�)�ce��2�R	Bb+��.�WwO�$����I��p9�(۞�)�d��x('����*��Z���R��cK��-a��J��m����� >��(õ1��"�~�S4	lV����U)꜂��5��E/���C^TYׂM�&��+��Qw�^�@�T\��/� ��HO��&�̡�G�}�bv=�gv�-�);/}�ѩ	��z^[2tgT��|{�W4x"���8� �M&|�}�;��>g�Ph��&S���Q�rևkp�H`�L�ĴYC�����Ti�ƪ�٬Sو��_趫��Ӷ���ˊS��!Gɫ'q8�����V��޶�V��L�`n��i2�i/���MW����w�W�~���o�I�_1b
�0|8�mE�Chw�QA�s4rZ�_BY�F����LZ�(��l<R��'������e�j����᎝������C�?���k��5����6������,]�(8����1|W���ICa�b`��x�EZQQ���k�l<QWX%�r&̊�>��!2��qN�k�EsqS���ٿ`yk/ۻ�ݸ�1�m�Ю�.�cO����}Zg�:l��1z`0�P��Y���z� :(D��J�����n�p��{�eJ{H"�::��AL�;���S��{ˮ���c�9kT5�4���������zvB<IF��կ?ǧ�����Ǟk�.,��+��'���Y��ie򕰲WZ?#�B�<0�u�B�jb�v���9F6�ɸ8<�Yo�%�̝��Y�0��n���Vp��_���L�)�\�n���"-*�}��	,�^xI@�-�&��p�����@��
�b�߇D�4�Lb	s��ׇܹ�'$�Oz��=4��>�>��a�v��e؝�t%������{^PD��S+�>;�����W�^��F;���- <��U:_����y$[؎����bY�.1���Xְ;x��&�om�V��*	�s�8e����[?�[��J��!�o�]�p!�C����{�0IM(x�\��a��<~���B�we0�N2P�|t���7T^r@�9]�ϞV�	���k�F�G�-��8����r4��^qJS����&oQ��k���K�3^�6��r����%<	��H�?5�,��8&\�8�aH��A��lD�9[&��xN22���c��n�4���?-R��L7�=��i�bdo�ҿA`ET��>W�匼d��Jc�EK�6��/�FV/�:�C�@6-���8�\�v����8qq|e�U(vd����f����ɾ�􉮄\�eI�P��i��h$ �Z����|��l�H5W���ؤ+�S��{����3�lI/o���X���4�������E�7�"լO?�.��������$� �-��i{�7����0��)�����u�ak���4�آ�v���Ex���w���?|�&I��VVx<׺��O�
��9L�Q�' �ԓ�{^)�ev$̦�@���ߊ���7&�E�����2<��s̲-&n߬%)^�܈���0�G�`�Y��Rn�vC���N&���>���1���wi���wU_i�~��E�����=�-uA�y�!�AP����� ��5��F�Vk�#����(��HvL� �ѣ,Y)�|7�ȵ[�#�V�l�-@�V&I_�Яa�1��G=~}V4�z'm�ָXW���L��g�0�Hǵf�w��MW�7So>'�oa�����<��O��"wȨ�ӕ`rl�\Ք�ݬ<L;ƫ�d�T&��\�װ<����z̎�`�1��{�S�`�[��b��P��l���Ԝ>ճX��];�
��U�VH9�sG��0�� �궔�7@�H��
�R4�VA�b��7�@�}�T��50���-H��Co7�/Y���m�Z6���!��.1Q%+�,����K���_�hEz�Ng�V�̍�W�?[dSY���-ߨ��/�2�ْ3�Q>΁�]�s!�$���f��CbA]0Q�/2�O�Y��ikrtN��LBA�%���?A��
��ƀ��N<�p5y���+I���( 
+<E#Aj�48�Eٚ��G4h�Lj�{P�ל+OX=�')q'���&�e�=�+�7Z������
Ie_ꝛ�ݜ��ub�w#߬x$	a��ˀ�.�j�=^��ƺ1J�O��K����~����o�_�e�W��s�����;�Wʨdģ���N����99����;��Q��y���,�@[]I@mO�b[��ߪ�ۇq]�[�@l ���hjs~o[o�|��T/��9G�����+d�R�=��~���h&%4i�%]StHj\u2��i���$���������(�UC����ʄ�Ƿ�l�eu�U['9����Ё�@&$��"HUF�F�~���ގ�TX��G��'LG���a�lZ4���F�v=iջ��CRVR��p8isPw�c�~�׻X`����M���K-
��$��⓵��/�®�\O�g�m��M7���U�����d���D
G��t���CM�c)g�|kJq��ޘ������|�-c4[V�ug����r���q?a�jwY�\�^���MYr2�gܻ#3��>�5R��-��	�94ᚈ�U�ktK�0�&T;�]�;��I�M���1�d~ȃl{�ɕD�w��f�@�<��iK�����9�I �d�K�Z_�rM�0�rE�Ve��M�Q�r���I�SK�j�Y�l������h�EwF����-馒,�"'�յW�s����Qtu�k��4�b�]��eǪ|_?
j�1��y�e�v��qJvf�+Ex��N�ڲ� ��V(q���;�:i����@Ѧ�Ҩ1�dP�wu,��a��ۣ+�Y?\�a\pҸ0ǡ����=#'iM��F�E:�&ǐ�o��P*P��ʽ�/���F��T��w�X�JZ�guh�M8�ӱ������|���Z�����u�W�3�!Я:��x����A�������I��z�_��f�oh��P���ԛ�VN@��=�<�e�1�^ѰR��1	���@u$x�q*������Q*����v�U/Sڞ��#;j����:���4��ߘ��L���������_�rī8�Ԍ�d�ӹ�z�\��UT��{��
���q��v'�&�����v���Ac\��nB���ϭ�L��i���ʛ
�n��V5��胎R0Oy��&���͘"�T�����!�_�#x����7U^t{����<��7�����w֓J^�s�M6��I՟�'��ݴd�bo�DC�\ԟ�4���}Y��C�>p���e�bHӔ�J`�e �����38���3@e��b��/Ҝ��ܥ��
՚�6�ɿEb?��ۆ�l}��1�����U�ԉ��)����+i�;����*i�0�@~��ve���]sN僕�[�������,�<C��~.w�R9����t���Q*R�-��1V�Pr���PW���a� �Tl�Y��q4���q5y5f�<X���Q/����O9aә��Dk@r݋U	�tï"�"�ԱO��a/�P"!
S���)�Q89�A-'���Gr�ԚG:�!�k�K�>ƺ�E<"_W�y�q������偡Q�e�SA���s�~;��_A�ʖ��sBh�uЗ�,�VFZ�;{'߱�<�Jfu���-'�> �@!>��0l��AM'D�5��a �Vb��A��:�UH��rw]0�j������4iCJA��zg��젦�	e1ϖsy�R��H��$2��ON���X�#�FF����C�`��k%!���n�w
{������`��L>"4�tO��(�J
E?�Q-Z%K�6� :���+��`����ĭ������>�Yr�hFrA.��	�͵�PC�����v��*��:v8��78��QX�%�ˆ�Xt<) 'J��	t�&�ۋ��e�
��m��s���t�o�Q4D��(�!��9�S��r�Y �^C���r��7��\�hV��ǟȑ)p���}��W�WП�#�
0��X6Naڵ�����~@����*�j����<c��nh>'_Z�վ�WB8PV�ʲkDE�^�_I�q��Ǘ�K┵���St�+Q�,�K��M�����`�R�@��W�W��-���ӌ�`�(c{N��p�0C�v^��`���ߚx����������x���#!�`���\�5��[fMq���EW�ҲG���}X��@c��8�`L�X�~MH��}�kU�/Ϋ����pӖd������Y8�����xx�s��cms:i�}��/��\�#���,�_���q ���=|��mq�S�H���,+ډ#��	8��Oyo��U�i�o��Nݥ�+�C՛w��]G�&_��䖐!�pG���ca�I���C	�PpqeR]��|�.i��K���j~��7��#���t�����A<�a�3v!�*$Y�h���`���≔����C����A�] �{ c��9��)���H�Dq3&T�k�5P�L���8���(�*nݽ�&q:<��4ۉ�f�Nt\��"%���m?q�ԬW����&C�c�r�W�T����N�Ù)�i_J0<g�����Ih'Hjj�����p��ӳ4d�a�����W�W�k��(Z1�[�*X���$ks)1�'�	+5xɃ�k��2D���m����2�yz�ǟ�@M�yM�5�Cz��0�C	�D��Mv�%�:���7����}���f�����C䜨��.m%��&?ȼ!9��߽��'F��.5����
��+�2�dr[m�0���}>�߀&se_��O�J X�K����ok�T.� ��_>Ztd8_�l}�/�i�e��L�c���g_���P���8�ՙ��5��d	�n=KZk{�Jˀі�L�e���x.�Q�O}'4�9~G� ��}�{���5�Q��L���-g���ǫ���j�n��!3�[p{F ]�Ww�(xCd͆S��#��ڂ/2�� ����1d�ExX���(��6�\�`��sR�V̀�l�i�MI���uJ?�Axa�k�*j": �� ±�K��a�ҁ��¡�<��D�V�yG�H��%)��n��m���y$���7�i#��F����|��F����Q���S��cF�#�׿�,'��SA��2�Bh\>�����~�x����6�1Fcg�.�'�������&��[��|�a��QY�穉�X0�?<� �#^m5k_,���2V�:�LJ�U5��) �X'꘯�Yv�A�S����}<b���ss���\��䂡�K���3���jK/�mŁ�G�ԉ�S���zJ�f;�O�9A��%g֘�3��5Jy-��U�Ne�$��R����q�c/����-y*��6�W����n����D9ʵ~������Pn��F����*�!a{�:8�G�^s4�WdC�
�y�v��ؔ%��X�d�3��[�Qec�ݵ囫^��Ӻ�ǒ%FT�OOzj*R6`U<��y�3�2���뭦rq�055����(
b�)��y��2j��	J@�g�*���Ve��O��ͣ+���Qޠ�qx2<����.^D�~5s�$=sP���J)�c����;��O4k�*���<j�V3z��_�t�3J�؍��/B���\��oW��V�Q �D4"�]��M=���c�~�q����&�L$����/!Q���V(<D�p�*� �"��Z:�}HiW]�n����U�~�C�BL0�~�{O{^؀5�L­.e��)�$Ћh�D��铰���tE�������d���:gV#���1�������7	�~!��?Ќ��	���`�a��9����%���z�|�'*�����ߺ
UD��$
[J��"E��-��KPfD��QI⊯^���y���-��� �ꡕrOq�_d����Ns��������0�A.5Jfc����gx�0~"G�|��ӣ�].V��#�Un�*�������3���*A�l�n���9�����ߚ��=��b�i�#iP`�G�(����?�b��x�L��DPV�^ ���mpl�����"���+���hw�%�T�D��A�	�qz@������7�١g_ܬe6���~�c9�6x��f��ɖR"��Wz�� 徒�0����,/5t�!_&1]�X&q!���eE�h&�W�j}��w񏼓G����7��y˨� �@i@�O#��?��&�]�E�������b��B���[ۉQU�~�\ֶ{U&��Z[
�r��C<0L��K:||(ndǽ�]�����r_3�O����E��E"	�d���q�/i�PX+�9󉻹�h*M�T*[TnPK:M�1�5'��,�&F�y��hm#�</\�Ov�u/�1w	�C:#pe��g���6p04���[*�qa��)�V � �m�C�,�fe�~.�ܳ�A�����j����a�׽jR�� ��Ω�!�gp�'�o���un�KANIu���	6���9"��@o�+��-C���_��K���(���i�*JE^g+ɟ��P|ѹ3�tEuԈ��ib����):�I�� �����o+E!��s��;/!/�XO��f�3G���a7�k�y �sl[Ð2�#�_������/�����_��:�sfD�ë���U2fW�H�p��'()�r��2��^�\�,-�	��V��c��K�݁0:c;X���kԨ���`����1���Q�����;�x��ctM>ڒ�w7�����X�Z�#oj	���2w�}������A�k��O3�^���v,�K��6��F&Şɨ�o>=/W��Z�rG�{6�h��͕y��^zC0Nj�9�F*��@�]U�P���t��[6��l�m~�u�Ӭ&���w�}�T��g6s��CW���}��,����*݂�A8����g^���a����wִ��	����.���po��:(���#��}�⮐D���[�<�o?w{i̱ N�:@Y�2m1����=|7DV���P�Ca�(��_�9�z�^s��$׷m�h&���Oe�P�ݚcjBd thϏ��D/����C�Ƴj�$'b&��Z���t��%���J/�}�U[�	�M�Vr���&{�*����^r����h�V>���m�
'�;w'ۆm>�QD/j�G���h��
Gߋ��+��4�(�˱I#�o��!+�p�x#"�/����G�d��Ҭ�����3�3*�C9,
y�ds۲3Vd+	K�N�VO��3���t��Ż�H�[8yCb_'�6�FCy�[c9�[�;��:aвy��1�W��ϳ]��-J��.݈�Eـ#��� �X1�9���W���nY�`�o��u� ?�&#����pņ�d"4Z��Ë��Z�'����-��Tp���rᲩ��)b!
�qj�k��fC� ��5X_�%Vb����A��P��P:���,(�}j����S	�S�jGxX^�)H9���_�F*&�i+��7Q�4��ڊ��������Bt��uXo��_�#�n�7C��lV���+�CڶPqw���H@?��I��p���+�i�D*(}jⅠR�y2�yB���Ok̯���ҟsۥ��56g�RQ�Wf�L3*������mR+N�.*S*�8��ԺTn-�%bW�rl�خ&=�`CM�Y_��,yt�����/��Y�Y��F[L�9�Wx�c��S�b�+��`��H�P�E�o��3�.j��<q��zs���`�cw�� Q��6���mL�֘u�"/0���ӷ����RY��S"���J��N�@*��;����]���б\[�>�yo���p���U6q���P�e�\E��a�h��0ڇ�`X�M�ж�-��]:(��M(�N�k��Y�d䂺@��EU'cDN�Ý���w\r�7:�N��;1�����P�h��\i;�����E�XxU �e_���Y4D�O/��?����r��ɮ[�q����PݟX�B&ш@��_`�Ф�� ����(���R�]� ��/�zy�6�w��բn��iڭj�|�Ni#L� 3��	3G(9,�4�><Y-�ʆ6���}K��[2��_�Z�0��"a��]XY�I����g��'�7]�jrj�Ov�`|i&z@cK��F�r_=zi���b4���Z�E��cB�@���QŲ�F[��ǜ�^ O��Ԋ�&O���Rh�s%H\!��8�@F	啯���l2�1�������9u�0%8�&�IrZȅs&a���,(�p��I��7K!�:�\l��y��ż��x?�������b�>	��?�/�l�M0�=D�5Xu��;��B\�>Pl���MK��\��ONn�l٦��1�$\�V*K�L'�2��F����O��s�־��01<�*|�4�\V�QO�?�n�M�Lty!E��~(��sDLVf�e��.$!�΂(wI���x͒� ����N�Y���L-3�* ��x��h�fw�I�:`�e� ���S��C�j�5�	}�3���7^m(�-2�&"�������"�*�Ҽ��∵�J���ګ�O�|"cw�	��4OǶ�,��Y�z���b���'&]�5+��G�5����첅�c�s "CԽ�G���Uf�O��m�$�� ������a4F��:�r?	Jb�UMC���\�燉Gk�x�_��>]�|��Wp>]��ى_�<n�K�5soP�\G����6�������_��{�Z��q��9w��+sT$R��	?�S�K���q4�7�<n>Fլ��޼L�I"�~�<�_���BWǇC�+���B0C���|����)@>D�	�� �H#57����T�	��7!(�j��0��X���`��?��uiq�Hև�L]L\W>"���_�t�>�I+����d@���������A���yWR T%�[
�`~�>��+�
�|�(���?�n��wi�\��Q��oO�ǲ��~;�xf�Z�Uj��aIg��z�?fMK���%`��T�~�m�Āc*ˡE��u�kw_y��#�g��
�L��:1�`+<<�6����&5|��=�A8d�Ƭ4��؅Vx��̢�\�7�� �p�	���^��*�y��?x#r�	ǐ����g��%r��ԐT�B[�Hj\�{��>⡉����}�U��uc��P/���'�U�2(�T=3VOL�u�a���z���pm������ܿ'P����S����eZF�2��p��!YkĊ�y���{m�a^�c�S���'�ln�e�'���[x�� h`�t�h�E-�|�DB����+uTN�K���s-����8��c{��j�S�;ҝ�W�g�I 8�݁N�v|8H,
)	�Б�<7������r��L/��6�)9|pvl�]c_;ͫǘ�J���Gn��~&���lGq�f���b\rP:�I�OU�7N���ǒ�p���T�>ʎ�#D�(�D�i;&�W4�e���`�ۼl�^����B�N,@6�t,��Q�j�;ł��b@��O����`ÏV}���!��ʐ��1[ZN�CZ!�M(�?V����G�ˉLz>�xy��J��e�5}%@t>9?�B����GJbv2_�e����;ֻqU(�9�� ���Q�#�6N
��PY�;:��dج��2�L���I3��'������
���>ac�
�(���Pu������$⏂;�%^sA�S����6����b���3�k��_*���f˭��5y����j~Φ,��K�%˧�G�d�=�u��`�6��,.��A��i�|/�V�Κ�|�ܾ��߻'i/��}�y5�yr����}X��&�$]a��K��8�R�,Z/���|�{�\ L���C����:Z�mZ���G��Pο�}�̛;�2j�������}ԓ����֠u�̚B�^@��bp�G��-��������-uƌ�zx�\��u6dA��fz�s�R�@�� �h�O�\��K��[�%Ϸm����މYşg�T�Z}��"��T�*���؀�k$3������'���k��
�}X�
CS�������{4�a��8�����gƲ����|�>r��Rj�E�B��@ �Xt�WH��Il?t@�$|6�����o��>��5��/YV6�BnN���]�+S_��R@�˃�羇G�TF��ņ\y�ݰ�>a����p
��nݢ�5s��1�-^V]����?���	��OLf���y�mf����l�ߑ�v4�l�Z���L�e��䨁$��	!��M�}:_�T�H'Z.���;�����b�`u�"?=��r��ZJ��8=~>��+��Ǜ��C����9"<�3�����o���γ��%�{���C�_gE}�9��^�m���X$}HsY�*��X3T��i>C%�r����}4�ӳ���eN��{����M��\���L35Ỳ]�;FT 7L�S�VFe�}��k��q;�bo�3�d s6m$\*�ݰ_�����ﱃ"�T����$����&�u���s��K��Y`�yqZW�I���snlV�Q���%t9��|��g�]��H���IH�,:�#��d�ā�
4�k�7_��
}qn���|��i�Y��@�P�Y��l���⍌�JeW�坎���Y��$M����wu<���Qi����ԊtDgmȶx�d��v!���ź��tucO��?f�r2���!�#+���-��	�r���{�u������* �W=�bd�q����x�C���Z�]�a72��Z(Y �¿���Xkެ�/b�u��%��S#��5pD��?�
��r���/C�c����s����b�)���P����#���E��$�b��z�B���(��Ç�,�T�!ZZq?;+��-��]������3�ޏ�:ӡ*/�)blE\��y%_5`GY$���*ϮSZt?O�����S�J���j�I�^���y)���Ɇ��LP��oU�͚A<����;��6(E;��ۧ��y�w�EM��X�����(�ЅW�����ź�`]?��������q���(w��3nơ�Y�ֶ,�F�����ݻ<EG���w��!���P�?��_�k�~�1�c#��?^����ޏh'N?�E�_��s�?E4���෉y�G�Գ�V;�]V��7A\Q8���x�֔9xhD�˚�]{n��Z?���f?6ϸ�lr�bE�U�G%��g#qoHc��D�]���c!�`�
��K�5\��[�:�ُ�v�]R�����MrIZ�������F��F�p2�����5*+Yg�X���,���%w��\���=�wOM�ɟ���y�z_�KE�����[�x 1l��>��g���f��� �[����H	�H�vjU\�4�E�)��t|��d�7���)Eʵ�/�Ҟ�Wd��FHvf��(���g�
� ����@C��q�
�$0���Hr�����߼�"P8�mV�yl�4��J �>�F����D~*SX�aM��c,���k�3T	~b�7YRwMeߺn40G.�6f.�P�c,o(����`ֲ*�9e�>I�K.6��+�n�*�x����#b?B�1�#Rt�NJ�����kl�A��x�pڪg��Ob�ޥ�*�WHk��LfS{��潔F�����Ѻ��%\���(:�@ih!$k�5�W��eM�=�s�ȝ�H_�&�Rd(��H��:`C¾����f@�M�O3H����l>pʡS{�p]�g�7D�Y���"�9H��C�2��=������db2�d��+��6KS�o������Wty��%>��\��0�a�xB�'��%��N+�*6mI#��T�*`&[Y���� �m�p���O���!��6UM������0�����O�u�s�F���/�w��4-���PZ�W�z|>\�$H�����Q��
���<�x͎�O��V����7I8]G	jZ���g�:պ�I��h���VM5�=�KtI�N�>��\�B�	.���i@P�9����+���JNB�� ��|�Ж�%y�4��v
�K � �v�3�L�&m^$d�k���p}<z�qVsH�E�)A?��F?G�lh�Xb����9���ƿ�3�c�5�ZV�8��G_O��ié^���F ��f�OD
&_�Ӣ�����?��[z3QpR
�@C�`��a�wQY!O���wI��CaR���r�@�t��̱�*�T۬ͫ
�%Jr�� z�\G!��cw�7ѢR����@��7D�f����k�����.Ps�3Y�dmăv�M��B���X������T#�N	���W�K(�LR8w���[��l�|��Q��<���N�(�"{���6q�Q^�Yk�YK����3	�#:6-�	:�)C�읅�a]Rf�iE����K߂ܖ�5���F�=#ִ`�

v[��`FTw��d��G���
1q�pa�gk��s�t�T�'�=�ر�0��	?�8��y�.oԛ��I�I�J�A*��XBˊ�4=�G�X�7��-�kSZ�UIVӫX��wJ��	'���8M��cu4��X�2w�h��HPG̮�9N(�蓗�{�ܫ�w�%tn�ڔ-ؔ�W���d���̢+Q�%?/�1:�zġW��%}Qwx�E)f_o�`g�����/�e�Ɋ�*Y��^<v�=��m%��A,��EV^JEzi�^z~��O�4�2OXM�j�¢�pU�A|G(w�z�)C+��r��n�_�I�wV�3G�"o��Ȱ��=*����a,A�C1�f���cCZ���cw .Sȿ���f\�HC%,i�P7�P�c��X˔p��_�Jw�Ic��~q=�x��.?�C\o,^���l��aU��I���w�{(;m��
�ǣ��+؇I�Jl�:(��}��S��CI'������G����6���SB�m~��0��UncY��!�	|��T2-��[���+ݲD�٢�!*]��Å���+*�u�K;/Z[y����̲�I+Va֮�)�@�Z`V։��6h�J�3/�I���Q�'( <��v�]�*��Qi��ڄQՔvP?��(E�PȀ�h��#��̛��&������ݜ>�*��`�Q����Tԭ��A�P0o����Vy�&6b	�R�,r��1�)�o� �=�r���/d�A5(��$4u�������a���/���^����\��߫��W�"a�RSJ���(�:HJⅉ�ߦ�"���db����6L���
RIp����0^��P�T*I��0C�BzFH�5]sɄ�2W\͓<R?A��{����
�ٺI.��XS��'}���n���.Q-�+j8W�,�|/���]1�JK=��֙���#�� q��:
x1�eR��~ޢ =n���X.��䉻 �Ž3c��7�ű��O�vܷbQ��/�	�J��%g�j΄��C@���-�ah>���6�bd>ۇq��VI���GR$@qһo^�ᆴ��椒�����$�"����_���v�8ɯ�h<���G1��7pѪu:Hau��HiK��Ă��� �1�1Z��\�>�&�votV�]_��W2�}�AO�w}Ք�v���+�-hw#�g�N�(W/��$|�e�/���!�rJ�����.���?	r|#Lr�(��lá�d�����Ľ��j���|3�B`�eH#���F�Z�̘@-��/�������y
G�#�ʩɢ �~%�b�Rl�N8� ������(a���Rvͽ�vr�*�&P9v�<��� ���x��F`V��35�*lߘ���͒n�I���T���qkr<�}�҄\����"�%������0�I���	��?�.D��_EÙX��rM���6��J�T�N&6���/��#�!X���>��Y��!�o����_{�[��m�7�̣a�����~t��]����s������M}j��4`�c*ZC%@��c�(�.�6���mN-Y�.�ň^� c !�0)���3��L��py��ëMV*/=Ԧ5�>Rnc��9!�E����2rü|��t,����%��̲nB��k�  �9.d���y�������uR������9������;��^j�I��i��8�CN��J��.�3ھ�a[{'^ F4m�z�QZ�{�A:�%�������P����i�_\�q��kr�M�i�Ӣ�1-5@G�z�ԗ����^�dˎ`\x�%��q�(7Q���F_C|�qZ
`�K�s�[��I?�X��^�z��p9`�����
`̝�Ӱd��"Vv���GVU������n����p���L)�g��!\:O�/D@��l��E��l�&��za��i������j��?k�Aa��P�vH �fe�5����fڥ�$�:8S�r����"�!;�b�e5$l����6��+#��<�Zh�)�
�}��)�����8ᥱ�W�ˎ��+��Z�~@xi`�B큗.�7��M�,���0��D=�V�GZ�R(�\w�\⛗>��9���b=\�{ X��iE�Kڇ��Q�&�w#D����x�y�6��DsN@J���@iA�	�_4 �7=ݿ�vk(�ه5%r�N`�0�#f{����/��u�k�����[��"o��'��X9��{@�#���|sq�����hHr�7��M �t��Y�oȣ��X$�	2���JRM���!݅�*Vc�结^^���ɝMw��nT��8uS�є��9�`��Z��8.A���xŬ��~Gw���qU�:gT���>��C�j�~\dѠ��@ *�Ɣ�c��ZA\ 	�
�!�O�!��� �x�ekْ��S:��_iSm�����Y�A؊\������~o��V���QUڗ��[�%}{��^����s e
鄵�'����X4�W3�!�oc�:�5<�i�_d�%~\� �
}�.��y�ii_Mp��$-H������c��F�)Gk�A�����+b��Yꤛ�\E?��w�,7ED�QoSj����@�h��J����#��7��=z���s�����I�t`z���\��B�_=�j���y
�ά�j���Yf��8�!Nj?�꤃M��s�`�lm�l,�/j�F�6G�Uk&��\a�u��^��y����nK�@J�[I )�?��ޤ �~�����4�[j{�_��6�i\�<)�fO2|肑�=!~iN����(�S���#S�v�d*��o�LVi�IY���yŶ��j�_Θ8G�k��2��h<�A�����u,��0�≧����lb��s%ŬFt���R�94h)�B�pj|nX��U��Yl���1�{�	ɼ u�`C�fs�@�?��koy���մВ��c\>�nU2�u�$za\�7������ȗ���>��K����lR�\w���@�NK��ӄAu)"�P�aP|8��
��r��p����Ƥ�|a��X�>�s&׳:27~�5�ʌ"�!ŷo&�'6�5A��5�����ϙĴ������=l7r���|u'���\k���/g���]�-V�2���ٍ��������xa��h� ���e״^�<S�����)��n*Gz���'�y��D��wK�<%�`���R��;8+N
��p��j&/��f�o���	�ȥ��Y����grN��=���`�w�"�rqt���	
�����9V8�q��I�@f�w`5���� .�*�F�������,l�9G��:I��s?Q���e�i�;!1/���}��+q�
��Fھ�Wv�:�&g�v)��?UU�����mT��0�q��C�Ӳ��xj��^���%p���#��I�m;P�A;C�]^y�/]�`��a��Z5%��gg�. j�#��S�-(=y�<���M�����ujJ/@�e�_�s%/t�^���"2YԬ����%���|�����^��(�g��e?�$:2�oV0�\K��Ӟ֒:�{_䫽�MZr��)�H��*kC���7��\�I���ۈSM��v��=�͗%0��oh��(���<�BH��\�ˉ�i]U?~��#jJ��a	�&K������V�CIL�Mpqx=�f� (6)�s{��<�Ҋ�Ggm�L�Ļ�*�Lq7�؂�r��cdCj�����K=�Q���@+��$s����֪��:#	wSZ�+��qI��m>����l߹G��ae�' ��	���^n4�-�[��TP�������[����䠐P�b�����!�,��8z�G�Q�rq�LWg%�_���S���ԁ��GHb�	�,R�	��9��B2-�Q�g����HP(,���u8Q��"nX<Ȉ �3e�q�b�>1�x��ǀٓ�x1�+^e��}Ͻ/KًM����WlN寨�J���v��>�����`�Ӵ�@B~.1g��u뵖t�Cu C�4����@�gBnPS�ΫN^;�E`b6�"��8Vve�z����D��\cr/����pMř�#E����H�wh��BH	�|�w( &ixm���g��k��H�/u:İ����]��@�1ZhԎ��P^ڢ�szV7:���=�VQ�9���95�15#��^=Vm9&v[��sX��ZIf�~�ā�X�^#���;���)�i?�1�)
>�:�"�m��O��)L�V��4�fk!��͛�����f9"WGq�����)�<ڝ3:)!��a�h(��\�TaGP�Mb�,�����r�\�ꛂ�����m8km��U��^*H��@����kN&*���#*�JO|>�R��'�]X�ء���[�:Wd�5�6�F����5�X�n�Z]�1�$�͚Z$�S�R���/�`܆9Sr�l-��DC�\ ��|���Il쵃��$�>vuM��8w~p�W*��#`
8�
�T�1;��)��g8�?=V�=�f�j=�_�AnG�@��]�TA~�*D�d�YؑhU}5E�������Z��Q��{��h5׊t(�Br7�{�[���{��_=7�//��w��{,Ϗ�ܷ��s{�M�OI<�㣁pА�z��[gΑt��a!<{�3�X���!_�
5,b����F�����%{�AF����#k=��p��I�6�`��;Hc���H��-�$���f�g�+�:OD/� ��֬�M%�!/_Թ�/P�Ln"�ËĊ��%�q ���+�]w�o�3��aIp�C?���Mn�"��C/-v����u�0�L�@�w��R9I��1�)̌I�}ߎ�B�����=��Q�����ru3L�HZ��ye4��ȷ(�.�$��Q|�p{яS�ӌ���Wt��ǧ�U�c���π:Ԧ�g��ݤx��e�b��@WU�V��R( �K�>��t�m&�3�����|Ft9nH9��+^�x&Ş�Z�/ճD6}Y+j���ws+���T�ӄ�M��~�6=�@/��M�q�ʢ�����#-���3�x4`�xߟH�������KD�L5��!�H?�c��Ǣ�S�Ҝ��K��)�m� �� )��58��"�Ż�C�r,�ë�!k�CSW�L:��@�����3�gE�x��QL��1�ǌ����#��3yY�*v�\֯��?���PP}	�)�5=@��FIE��n���@����-g(�l�D�-0�2kq"���U�/&:N��b
��;�Hy�JR�^�_�L7�|e�f��������X�Y�H�)4��P���<����*D��s@�a��%v�P��)$>�tCά��?��ђ�L�V�#�Jk���9�)F�,�����������p�(��چZ<����EZt��6��	�Kr6�� �cY!���#ָ�[����K͗�!�f��󙖍��!�*���``,��c�m;?f����F�+!�_-4�B�3r��0���syυ-�g������/��
аm!;�0�P�$p��5ZrQ��W3׸2+$�Pc�9+��ݨ���^k鿡?S�.������@��2h�dYM���N4�~.�iId+O�_d�P����Y���ġ�dݡ��l����_�7e��u��w�y�F���2K��O����j��?�x���l>I�^.��k4��
���/���v���-�ђC��?�T6~��s�V��_��e�0x ��z�-�b��~����o�b��~R-�^�����a�Г7϶�%�`����ص��K�� �5}P	�[�NFL�7��Y�1BLl���`��ǀ�?$���N�9�bȒa��>fh�?5��ƲW}����2�H�W� #[��U��)K�|Tz圙P4����
���~��j���I�}Oh��G<*>��ى��X��2��GI�ה��C���rR��%2��s��U�qj�4�Ə���oe ����_Fmҳ �Vu�U�I�ر~L�Y3��M��_˯�~���I>�hm`,����?��@�b���4E����tI�K�
ѵu���zWu����;��uhD�OilI���w�&^�����X.�6�����<�Cȗa`?�Li�����T#�j�9�A3�p�;������֨�nۄ���	�4�(~�!٨O��fT�ې#�e�9�k�hĘ��S���GK�'kf�&�ҠyZ�\�������S��D�(���-������C��i�[e��9���� ��C��M�i�LK6�!�X���@���~)&Tef'���'X�ۉ�,��B�֚<G/%�ґ�2~�w��jY*�L�N���r�Z�������-~d8����}DZ��.L�~x�R!-K_��&/�����L"2�%��@x�y���o� �4���b����b��d<�j��i�.ږ���M�����^qk
�yzG���@̔��%��@�����ބ���F�(��apy���b�D^�B@�x�."�e@g0C��9Z��:\盜�Uyaj� HH��F;�5�KL��O�H��jr�-*-��;�����c�'�Z�FF���6�N� �*!w��8Qd��;��et��s���^����9�/�i��ѐ]ٖ{���hH����t�[��vӿ࢓4,�0��[`�=zC�p�R��N��0P�c; �Vk֒h�[���_�� ��?\Ԇ���lC^� vM�g�+�����/T�P^�[�	�1���������M�	�v0`�9��V�x���p
�,ʚ������#-:��	��\������o�Z݂O˨@=����ǉ��ƪ�J�(�HS��>�iF��'������>��F�^��l6��`�b6
Ä�!2[�@��C�J�ˀ�^{���'����og�׮�g�?�X�dFN��r/qkU�o8tNx�?D
�EV�ￄ�R��`�D�0̳���B�TkG�V�i���4H���W}����.�WdWI��ľ(P���?ý�zQ�t�����H��}�p��AZ����B�7��#m��ŕhX�� ������YGx��S�R��p|�B�R/�.��*��tM��BH�`N�s�d����E3�v�X��QSrX��b��QY�D�sjYq+�l(gv�W18͚���,�w��tf���0�Y`ˏ�^�9JeT��	Ţ��Zjt=x��L\a�4��6�2�Qs�\�5�va�z��He��:[�xpv�P@>�N���eo�2N�$��x7;\_$9���.�"0]T<_;j�R�0�?a��uX����S�Z� �����?��u��8�)�W���"^M��+����J8lC��ZQ�ޖ\W�4�>�åu����\���%D���yԂ��gS+�s4bg)���se\�^Z�m��.��g��f��7u ��_�d],�hMݱ���l�>�$?�йz�nʹ�A�R֡��~��f_on �O����>cܶ;��|J"�5���0e���������xY��VH���E��(J��͚�6�$63��[��;��iI������a�� ph�0M���!%~�>�w�a�w�س	,��QE��>��*�tVA2�.�NF��Xs)P�ՋC���XT���}�C�%P�1)B����,��v���E��x9NG�`5� m�3�kc�9��q{��z�5Y�l8��[�Y ��g����u��*}�^�����\�����D��!5:Ӭ9����;�ë>i�t�+!RW3����O��[DV�*D�w�.��}'Q�V�|^�l��-��=�"�WK�������̫Q��B�N1A"��%���iE�	{ĘY�Ӭ�K\���W4���b�D���J����(�E{���Z�;�CC�lh�Z4�c�y���Q��&(���m�&�v�[X]���y;+L�˶BsֺD��~�^W��x�;���X+u�?{�(��tyWPѽ�>V��I9?��Í�&=��h>e��z�����/sF�>f�	n�r�q9��/��vYk�]c/h�9�RNT�f�|'�u3�H�a�Cf>,���+�J�5����S�<��]��т��L9�q�2���j�B�.��1=p�Q����,�ܥ�Vz�Rl�W�D��������BlN�����U�6�6���'h��z�r���B��&�ܟ���,�^�*���!�'�V5�\�iV�"P�^q[�R��	�*�l]��sW#sG��/y�\3�oN��Ћ�Nv������H���B��u+�3�/�·����'T4/f�P�6X��G*�"���'#FIKWz�`F��0�|������X��i����K{��稾q���<m�S3 0d��w�R��H�ƃ�o,Zc�	"`P�A K�^���?R��E@h-%��2ye 1j�����7ʛ�ƨ��;����L	e�ڕV
Hv�y��AZ���� W���ԁ���4�RkXv�6;lt��<N���VJ����Ӌ�y0B4=Ι�Ae���@�6'��,��~��oQM1�X�D�,��g��6Nֻ#�|�B>��,�S������c��������H�1ڣ�3\���<��{��A��?�1f��uK cl�_��������>��A�QoȺww%N�����z'(M:3g�$ַQ;��-�w��ZWi*�l��C��L+�;��ퟷ���_�&?����Zد�=fc!"��Tp>��hN�S/����e�����k�V�,Q�)��a����m؍������]cL=v���O���d��Q�{�5NZf��<�2h�LεR��+����f��Xs\�q6>�3ʱ��ʏ4yh<gx�CW��,��3�5�X�H�i�S@�.��:������d2�s���~���Pk/�jʞ��#=��svT�})���fC+��]�5P�E��-�\���zP�)�y��k���]�eyr�,�ܔ��i�J��4ܲ`��
�%���l;^��E.fm<��\�8gfW�1���f�:4J��-��χ�%
$C��nb�Bm�[���g����P>��<��l��p��oyaZu@{��9nS�Z�1�?6Axn����>N9&�[<g�^�ai����~�l��+�$�Ҟ�:�{�|
V��شxq�sV�ITr����8~S1��3X�@���8r�-TX��M����sNG'@.��zH�W6�a� R��ܳWN�S�F�{�m4��a��M��IL��5U�~H����?��iB�A�K�o�U��ҹ�,��x'<�F;�����h���
l��?;��?��N���G&ǐ�>���؅9�?#�1i0u�"qm��ę���������濕�?8����3NMZgX��ֵO������هO�X��58.�F������	�?�\a�Ļ�>"H�ϵ�n�E����e�xDe*Bt%��B���_v���F�m�ɲ/�����*"E=rltJ�����U�ֹ�4b��e��s�}AB��V�s��bvO�NƘiA�n~Aއc�Uh�Qk=�	'C4 �-nϠm�H�&���k/9��芀�G6<T����^�)�<����]�����irl�k���ՙv�l��p�-"l1~y˥9!�@�����8~�HrIQ�����H t�g�V��⎆x%���œ�N�3x{[o���Q��C����_�ߕ uԕ�6�=�k��]�5�N��=J�y<���4�z������:bD�9?/���O�s��6�ʣ?�|��k��]�K�8�^'.!��3���t{M�|�<�D^g�%�,��(����c� U@>�S7������N�1��;�0�1Y��=i쎉�iԙ��ϱ��ދ���0sď���.�d��� =%���H_Σ.�j!���)��&����4�[�V]��o\�	C:��:tP&{'!���v,�^�p)���]b��8�͸���Dyf郩 ��C�3��\�)a�@"���,d
��;����7
�y2��\9P��5[�@�xZ\~:m��kOo�H�64��/�.1��V��	�
h�J׭6,-�a_�+HC(��w����y�*����#�5-m�V����-���m��n�F eP�Ԗy�}���g0*�靑����ί-��ԉ�］��x�;2� Fb�k�Ž�e�gr�=ù�x�e�O��-���ު�d �ȑ��+��IA�s:B&����f[�����k��1z�[J|$��ѝg�U��)9��6�����[\}pEGJ<��_�V��������xx�{����R�Ek�_kQd��`���J�:ћ�C�k�K�����v[e��"D��� ��E{�%�����I�߰6��?��W���ŀȇ�B_٦�Ȉ�}��B0�;��	�F�F����1*����N�!�-�_�`A�A;/@�4�=bv�?���D6y�Z�S�7|2��}M��A����n1��DL�@E �9؇���t\"P��E���$�z0<��k����_٨�B���y�1�0I�ɍb@#E 1T�Mo�`�2��@�	&���By���+P�r}�ue|W�F�
����"�y3u(+�֟�?9MBT���9��w�U�>𜩩����4�[�#r��1��P��W��C�6=C.�,�!���A#�Y�fUv��ٶB1������f>��"*T[����K9|V����[`痥���)��a�_ŠXF�oc�5Dj��I�_���ͽ�V���A NO���15	;�y�xx����P{`-��گ.fj��/6;?,�;}��7NvsG`}��sS��=y����G�J��T93�����{l�{����Z�K��rE��F=����;�*O���y=J����ܬ@��Tj�:(���*M��ö�r���*��E�^0jG�ˆ<ДL�Dtb�'zZ4TYm���>��}��������i�Hk@�ۈ���%T�/�fϙb�+�$�c��&Tq��e�f�<+�A�O�!��ə�f�X�=��a���s��l2Y @����������2�bӴ�����+ٿ�Q)�OBTH���[���������P����g��R��#�/Z��)mM?F(��$#�n�y�ic��q~��g][T&�
k���`8i��)v�E�����!�1���s��iI�HkjD�x8.;J�_eOk��EM��;�֕ivvһ�%&"y�XH nCl�J����Wo���W�\xX���:���� ��j�D)��rs!�ȍ⮗˕�qX���/p�JV�~�b-GH�����������n̯�ͭ'�Q*ُ;�w/j�	6NDA��:=K�=���&ő��3殷���9��A����R�[�%��`ȄA��']$�B3R�����N����S���ʒ!+!M���Į3��P�˾M41�ڙW��-B���wh���u^�W�Ǝv�nAI�6<P���쓟��h@�*��Z�L�=�0]�����y�?�^0{����M��Uo�����L����`Qp#���h�q�v��Sj�,�ۊ�7�{j4�ܶh;5��B\q+�8[��T�_�<7�/a3Fc����؀�m04�ad!OK��)4�8���Z�6l8�6����~5)�~�%}B��H���h�&\���.�?��
�;u��HS��2�u�L�#����c����8�@bD5�v�9���+y�ހ?��U1��4HV��.g48	����o�L�S�T�Ʃ��0W�+�cq��Jꦆ��zk�`�1�!��D��gmT��v�ʕ��5�+�i^���@���^�3��v��k����)<ǩ������Z��a\Zf��s�`ڑ_���٠��Ij�4��& o2�~��TM�������6�f����v�Ջ#�6�n��S�!��R�E	X�|7=ǥ���s�J��hP��M�)����ˏQ��uנ��4�U��� v�11��Ǻ�7�*<��5t�M�4��!�A��d��2���r����a�z1D'D
+��ن�f�0h������t����/�H�[�럑#a����X�e\�ɏ��ы�l7�`���l�����w�ʌ�Nz��>|�ajz��ll�¸�!z=+�ȥtjv'JGx�<FsW��{l?/}i��H��F�J<H���r�HsМ~vsD��*�������P�m�rK�o�%�a:}��h�Ɓ:S�S'�g5��9��y��
�'p�]�Z |�y!�n����h�C(��M�L���X'ldBى���񁐻+I��]�R�~�n�������1��&�B�}+a����i�ޏ��Aqr`=gӤ+#WC��o�ۃ"�.�%��g�\#��lި)⣈<�盀�\N]!�h������d�8�X~a��l~�g�#�;@���Sb`�Oǝ$��A�(�u���?ۣHk�>���2����JݐB/�7Ď�Pq����@��l	2���JЯQp�6�ٛ.��D`Į�1��K"j߷�(Ѡn�l��QL�]8��p�-N w���]`���6O��u(9?@�!*%���R��d�J	RzqG���nG����+_65��x�_�-ɢ��.���D��/Hز=7/�0pٴ���ց_�K�w7��9���8�잮j��K�o^Totym�׺������ \%��}�-��3�mҘJ�֢$z���y�V�3~;��E&�L.�ͮ�*�*zB$���y�L�q��m�W�+�����~��u$u
P?J���NZ��p:mt�����Ld����I7����v�W�C��_����{�����3VP����`j��n�h���脣�xϪ�EFI�%)Jv�hAQ��Y��SZy� ���98�������+�V�w����0`�7=Y�0���_iQjY��+���=�(A�{�~��t��+�����n3��]��Ɓt� �M}��8�K�z��5��]��{Js!ws�~/ �"�J6�8�Ĉ;�s?�b[�Y� )&�y�w��N�5Ϣ*���~��BB���d�u�`.p͞J�JL�{	-�e�M2|�E�2�_�
����α�����~�b$eE!>z�����A�1�2��Wʒo�%�T��������M�"���D�����m:\���LYF>��z�J}5#�<B�?�++
��O���N9�%<�\�)If�/.l$I�ԩ�5{��}p��R�e"��b�{N��Q�&���/�Ԟn�y�#��]��|
�\\���+�K;L=
���:���]�ۖG2 l��r�M=����L�`��EGM���� yY��5��n' �X�'� ��rn�3CG~n�=�U�	eW�f�	 �;8B�'���y�Γ�Z*��)0��~9�~������5�K�TL����n_�� ߻!g�6p�j���nO֬��*K4�i��0a�s�-��dO�U� �Yf�NXW��z�5��>����ibX�P�Tן��d��!��<�zM���y`�)��:��(*Δ���&x�Z����Z&!��m��RN��͜�k/4�dl��dq�������r�� (�8ܶ��d9l^�"�'o�˟W)N%�U�h�)7�Ʈ&���=P;�� �H}���lX��S�	�i�ݓ]\�,�ѡ�������6\���.���D��[�F/�z�x9���ɣ�j�L�똎�1�hv��7�G����J����a�{�	��ާs�u�/2���y���ژI��u���?+�3q��-<�rt�t�ړ,�Q�ks=�/^#M��l�X� _��|*aa1�k�ISs�v�w<3��3D���XG�S��
~b%�g��7s��}��Js���dy�B`�Q2^XoIԦV}zuiCV(D���w�2f�xϔJf�,0w6�ߏ�k��B�b�,�8E�N�;GWP�����A�9��4��r�}����]JtGಾ=��N��]�.\����m�8�
��m�=+��\q�V�8wT�=��n�s�9� ���O�@n�1+�c?%��dL����0��g@�*�)rQ�������'��������� R�R?�-p�3���C�މ�4#�զc�h�,���1o���4~eG�t��hcM�)����Sպ>����e�T}�+%���M���m��^=��,����:�i�˲��WD4j���_Au\[vB5]�����Ѕ�p��>!��z��*8�������#Z�y� '���,e�;t�������a7m�J�au'#	`ܰ�,�~�����֝ӽ��@	���q7�9�W�����^�F��S�(��v��d�xˠ�y�a`Ë ����sTS c�K�o������ן	2��yO%���2�(���q��LM�O5��n����RϦ�g�nh�������~ny���h�ߎ�j���
Ys� \>�J#|���T��P:'��Qt�������X
t����9���Ҧ��8��44c�n�Ws�����.IO����YØ�϶]�}V;����`"����O�8&W��Oݫv�XN��?+�����t :c<+��5����~��A�K�;��}-�'I��n�0�Q�o��_;��j��)z��*���H3�.iIv��� �Բ�%̘���u���x(}1����#�Bz�3½Wu��o�$d�b�v�K �$��d��H�� ]Jt�C��Zl2$�/��9icGz�Q��#���tI��|G4ʢߡ�Zf�Û�\�oe�9� .��;�J��U���	k����Y��>��Vj�2��y�ގ��bS�RM>�W9��5x���z/6N�\ ��/�踡���#4��?�[IS�P�R �6�"���{����D���V`�7*X��Z3�G��Uxo������Y".���ə���6��9���y1P��a�����ț�E�ZB�g�s�h��b��K�f�)��qo�g=Jn�ofteP$�� �w�����2�nvϣlGŉ^�n��t_�{�6,�,ἲ����j
Ilt��
;/��ǿ)XL�[،w��Ymۅ��g�04eF_�r���û�Bgk�/�h�N�X�����9,aRO~aǇVylR:�Ș=mH�̣j����'"/ءVQ\6-|A� �:�
Κ��6KP��ག	�"�13��&�����T�Ȍ�?���#^]�F؞�	�^�p�ߺ�K0�G���n6-�e����6�7�:U��v�'�'�twL�����E����y��_�x����Z����C�+Ŭ����SX�]�T�)� ��8n6`����"�Y�	�]$)�çE�)�+k�LS3���
\[�&˜y6�^`tήav���[Hٱ��T�p��,�	[Wb����%�U�ɸ������b�6F����&�����T�vL��	B.��`�����A�����|�q�����A�r�K-P^�p���7�4�y���o����ˢ�$�qZ֫˥�9ט<�(�|/Jk��ϖ)��:��7�+��,����F n�e��|<��1v7B�w�X_�S��<��T�//p�<NǊ҉�U��P�g��
������?��%���\5 ���׋4N���X��훭�ͯ�xU���2i��&�#�RT`h�r.Ej�mL�Q�.y��7��sP�F��0Ɏ�&�)�.�:����ԗ���vZc�ժ������99۫�e�h��D67IB��۸򜺿\>�
T
l�L"�v��mW�L��8<���
��!�I�����c�`��2�\���>�eV}Al
P�B�a���q~b\���-�-�T�&F��򡼔(qz�-��y���f0Bꃟ�u�m��+VM#A����	���7�@ ��O���./SX��Muxi�jbK9��q9��Ա-�Wq|xf�|�L	2�[H;bgx��%�5�����#"땄9O�]���<�V��4�6 �z�W���q�Rm>Cx{U3)p��:�!��㮿� [�M�.'��㦫`�>@ּCY`��^`��ڒf�É��j�E�+4��N�kL�����S�-Z�cR]hō�1��&��J�/��e��c0���AXz����_�8Y��8�ƶ��/6�yX��IT=,Ͻ�8�)�I���<�WL�TH����tw��h�$Jq�'a/����Ha��`���-'��-3�a@K���a��ş`t��5y(�O�[�����̃ �-�9��r��feB�g�w��N�,t��\҂P%���Y���&#~��Q�Mư�x!/L���iS;�$�sD~m�3 k6����~��ՍIs�ю$�v�U����$�-Ş?��J���ux8� ��o�|s�yS��?k�}`.�_�D�A���z�������+��Yz_Z��˥V��45ʏT
����dT��W�M�t��Aʝ�_��Dr|%��@灭��J�qv޼��W�P�c!,��8n�'-+�$Nh�&��������I-�6�{���*�6LL� �S�+���6���8B������i�{&ǻm��#7���^U��.��e�}T�}[B3Qkj����L`�<����I�lȇd�sԘ҈%wIt/�����#?U�Ϗ�C�.�~�W^�)�W�HOp�����O�4�P�˗u��/(©�2&�h�ܪS5��`�Ŷ'��%� Q�J�M[�yI�FULP�C�z�<<�>YX3*�cIۭ�������N �Yf�o֋�y�(�˧�5�P��a�'(��l)a�JgQ�2!�����}q%Q3���~�M�UȭTQ
�)��k�d�_�$����Q�B�;��<����q�B���04��z�O\���e]X��}��U�	�G�v��Bxaz���RIܱ��h�<ݗ����v�M��kRˍ�)Nu�}�
��)�s|���DJ�ܒu�"��ߦ��A.��Eю���iލI�d��ȧ���3��	!	�V+���Mj��V�
���G�te��Nc��\��L�GBt�(�^þ8��B�V�prxKa��{;�o�3�Z�p�/f`x�yκ�4�D`g�AY8.��~F� ���o��b�Y~٭!1g�*��L�`8>,\�@�eY����cE[�blI����uay��i�0m=�jo�+F��'�Y<�6$�(��������paXN�=�W�4�S�"�}���᳻u�����(���N��Wח$�$��Đ�'�r�>>dC�d�h�} ��d�\�0I����)<�7�g:u��!�������_�!�P��3LȲ�r���tErve��3�a���3$�&�(��e���)H?�US��Ewϩ�ȋ��f���e%�������g������ř�Yd�/���!��l�>5��I���$l���D	n��\�m�Gh� �A^_��W�[�z�M5�0��;��Q�����L��.�"��:���z��O��4q2��W���?h�_����'Z~��nCtq�Vd��*i��e��`fg�T���	ӕ��|�Y��K[��B&�\�<	i�&5���15�ج��h��,�uS��/�҄s�R�\=���q[av�C��
����J�X$�����&cZl��`��7|�b.�{�2w��M�:��HYn���9M�$�r�J�H[�׋�K�s��������>Ե�'�2���Eh����8�<xx�4�>l�5&T�PWmd��<*�fڞ� .��G��4�=/<�s��`�pQK++4|�f�N�37O�&4� M��1 �1�
��V��:Z�#?%�]>ÜJ-$۰Z�E��r�^9� �.����T������E4��w�� �v�B��t���`	.��������O�24�IXs�忏[%!T�i{�g��0����|��z����@h\���ZydU�H���I�Ke�Ơ;�K���9���	�*vF����h�"B$�Q[v"3j��q 7�LI
;��$��^d���3���iT9B%��ʮ����4��kN���a,��\��~���g,�]���Y�4g5V�%4e9��UZ�*��&���j������R�Z���4	п����d��ya]8T�g�ɾ�&�+�\*�Y�jϴ�_��8u-A�.V�A�mz%+�{ܺ1�Cg�����Ѕ���*��Z�lt�_S���O"9��&N�!>�>�驄�g��P�+ɠdB�Un��VIfi��[eriN�ؾ�|��Aa{�r�(o6�jO)/�ܓ�?�D�|�(.+|�ᶥ�g�kXS{���?�.�,�B�2���5�qHgBLRZ�j�V�y4��-�dhL�g�)0l��Xi�Bl<u��6�d����Z9y�K�if��J ���'�����$]��ޝŢ=&i�gN洠�]�9"KA/��u��oO��UNȹ\�O{FJ�%&5���s$���;j`ӷJ�_��Sn�� ���y���KU���w��i;=��0i��O���@�4�m�N]��^�:�GoLѮL��߁�v�nH�g;	$���n�*��&9�G8����y�!i��Ȑj���d�?�-g0�J+�,�0�DY��_���d~�:%TCw�C�b��.D������;�o�Z��`.��>c�$�Dt��c
tĖ�E#�$�YzcgǵǵU7��yN�͘�B�cL��8bdKz�H���¸\v�ζ��U��ҘL���3w\�a�Ih):��dS�^���&�
�⮶�������E/3M$u ��Z�en�l����9�������v�iø��R?�v��\H�B����N�0��|2m�d��� �R�zR3��G>a�.�FRZ��$��;Rt�K��D���H���IFj9&B�G{�v9r�m��}��U%;�W]F1h`�����7+��q=>�i㧻8�P��m|^����ɲ)%�3�����?8�-�
"�qW!U=?�6N宏]Ӹ�߈���,����iΨ~�<��5u�`����]͗�����gtyy�z��� ^|Q�8_�.A.~7�5SKx�v&W���	�"�z:��}[��ΗZ`�7��(bC���W�bn�bB��\guk��8�<0Ř}e�w�|t�:?X������t�@��d,����êCc��]��[�,] �׹�!���ė��WŹ�nk��|Ì���!��TV�._�o5C3a�{�eO����63:
6�	� 'A�/}�X�zh����VC������+����۸Q7$�gK$�3,��x��{5�x��H�2`ԧ5��]~q֟!ug�l�|�}6�rR?��ܔ�x�ρi��rЭ�H+̮��.��%<c�Z�=SQ������}ڭ�b_D��:�����B�]�ꕔ 	�$R�#"bݤ]�s��ѳ�i+	��'>O'7�&�'��/gy姖(�y ����]7�BX�R�	�7fVb[� 4XP��.^�-f��Bu�y��櫆��uL�C� }���XbI8]eEe/�ʒ��!�,�|4�Ȯa;n�&�-�8Ԍ�ne�hO����5[C�B
�望HU#c�ɩ����%c���-������e$hᶐ��Y�M�5�KMF�c'�;Ѽ�-�{����Ån��
�0oD�Է���"��%�K�~=
�E�!�%&@Vb_.�giJ��u<0_�PRMdq���U1L�AO��ڰ9�NO,g�9�2s�{<�浡N��7�g�r�Q���h*-�������C�!�^ǯ�5�Ǩ2�Q�37���U{7'���q 8D��b��G��ܩ�� �̤���|
��U=6o�����-��p��HIq�UJ��5]�,������q{Y�5�_b�1�u�
�ۢ3Ko4�>�욺���l�\�NX�\3���d�@���U1t��P־�:�x'f�Q���ni�۸�x��gc�0w��`��c;A��&�9�)��}�$��C�ϗ�l��+h����f��$��<5��u�()�p��b��c�b(h�谤����R��Qɚ��Wa�WM�r��b#���^��b|��6�N�"N�2�[�q�%����H��#� )����Z�&���1��2�9�~��`��K:p�^n1�&/��|����g����z�y��� G��u��,l"�G-�[k�i=�ke��ՈA!xLf{����k�GV��G�(Ӥ5������8�!����%�\�<�j��E���0�-�6_��ڥ�����O�fr[<;�)a�D�Ȼa��b���|�-K�-�.!��LJJ��O�,�������3�e�Ç;������4J'\���c�%7��z�>���b[��I����AWA���ɜ`������0��V���s�����=��R��������`aL3@�H��W��Yz>rD�rHNS<ڐ�`Xk��d�P�R'�M���%�ԋ�Z�>
;Uw_W�P��O�YG���vbu������ԩ,aȈ��i��C���;��!#�N�Mf�.����&�H�YePzqϣ��r��heQ�2��K%W���,���q��C]�����~Z��hG@v"O7j�B���ćD3�V|6����3�,���x4ܞ�]�0c����H�`��x�!T�R�;���N��c��)�.��R$U�c�):RM[sYF��}�(����r+"�HeOO����+QɃ#=�#zr�y��Iw�٭�VD�x�U��&Ϫԇ�V>��w�z־l"�]Ѯ>\�{۱��K�Tc��B�yIm�NҧB�D�C	�-��<�`{ؿxx�\���8)���]�ǫ�4u&��O$@/e��X���@��˂�O^��UU��ԫ�����U�'�gƜ8����ٿ�[)����,<��4k��U��^w�p��q㦨���1,G*��D�@�=i£��n�{g�����/�l+ԕ��mR���)cC�`��Ss�O������T��h���}��~��l�H��
��?<!vY��=�q�@A)��fŤ!���� ���c�����q�J[ο�n5p�u��o�S��B:Vb#)�m��~���J���������E�PE���؟�4-i+�}K���,���=Ai�5���ߥu!�#vOÄ%B���k<�x�
[���1�i 5�U8$�#�I��R���*CPg%U��n�`-oh�K6�!e�g.����I�un.$��Ĥ����/b�ʑq��ø��j>��z1yk��r���|��#�G���j������ŦV��?�y�j&��+�^�f�YL�ؼ����&-���R�6��TC.?��iǃ]�i����_j�HH���l����r������槊y�k���V���&pWV^�D���p�;��R���2�9�=]�)I���\M^��"	Ӱ�&�o�-V�D�/��O�[�R�xA �Y7�q{u5��c:�U�=�=�O~�WR� �FX�P���>���i"�$��=u�:��V��U�Љo�N����0�Gj������7��y/Dg,ŧܮ��H���ƨAn���D��.��rX��4�^o�v@Ҳ�i�\t޸���YG�bK�z�/L4���u�98��w��Z�������ݎ�Ȼ�R����i��R{�
L���&ͧ�G>I���~�%Qs��	�wx�ֱr���7�H̋��Nz�T�C���Mы~qc�9/�-����6rF�������,��J̨�AT���m�Lg[c�lJ��i^����`b�k-�\;��0���%
��&��!��7ܯo��x�j3��q�5��D�����.t&���TC�~U%x�"����
�U]#��E����é�`E�$!�m>�E�����gAU/��O-�"��Z�p�{��h�v�IM�}�Έ($���s�9D*v]Wtߜ㕾�f����ʍ�A��Z~9�d�T#-�f��@����	0r[��,c��yKW(�x~�l�T��@٬0���M��(������TO^�iR,��jc�r�����Y�d�1q���s!�Z4��#F�`s����.S���J�⡤(	�P�ڛj@���V����2 M`���4�z�6S�j0�럹)^�������8F�D��O]aI�}Rf�Mk���E���^������jwu�����h;�K���z�3k5�?�Q%����f�''HJL!=Ƀt���/���zpZh<�敔���	��s����1*&����@�j-'dT�Ϩ�!�Rz��Ku(V�`-�5�2�y��MC����m��x�Ş��7�JGO��i_Q���識��׌�=(��8�:�Zi).�=��mk��t��-�'~��/[Ł�����*@��y�8Wg�Q��S���$�;d y�%���2Q�Z��3[�Ļ�H�rW�^�d$�_n>�us��r����"ܠ��!l���h�N������Z��2W�ا��NZ`J�/���
��Åj?���˕��\VtW�`�+����z(W�K�S�F��	=煼g{��6�.	��I�T/U!��N�B���*��2����T�v��M|>Ex�0�n
G>�� 2,vj�z���H���q$���h����ˢBm8
�Jhk�����j[���R�$�Ӫ�xLP(�nU`�Z>0�B=2)��(�(����3����I�ADE^T��T2�[:x�
'q݈8�g�C�C��qh�x@�T�߃
�wkqu3*�h.��on?�&� ����]y�g!�`�{
4{�G\~,�oU�gd?n8 ���d�U���;E|����Lw�R�%V�x�!��3����8>�TD��p���rT��{����0΋Y�u;'� �[6]���qw�	l˔��b��_�պӒ�3Ҷ����A�[EP?�������P@NL@���P��]��������Hڲy+��ۺ�K>xo�ԧo7�Aj���e�?FM����~y{<��%��\��"�\\�yo�DT���Oq��s0��I�͑J��L�1q� ,Z��p�W�=^*�ޞk����S�����6�:ߛ�pR�Ä��]Ͻ��R��$�7���O*���)
d�X%Z��	�	Z��E�����SK�j*�Q.%�JҎ����m0�A�W�t�&��+Lc">��凉5%�聸����}�\*|0�`ߊ��� lE>E(�D������>�n� [.�7�鞉��`����Q�~u���\�5v����