//Legal Notice: (C)2008 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module build_id (
                  // inputs:
                   csi_clock_clk,
                   csi_clock_reset,

                  // outputs:
                   avs_s0_readdata
                )
;

  output  [ 31: 0] avs_s0_readdata;
  input            csi_clock_clk;
  input            csi_clock_reset;

  wire    [ 31: 0] avs_s0_readdata;
  my_build_id the_my_build_id
    (
      .avs_s0_readdata (avs_s0_readdata),
      .csi_clock_clk   (csi_clock_clk),
      .csi_clock_reset (csi_clock_reset)
    );


endmodule

