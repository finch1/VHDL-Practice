-- nios.vhd

-- Generated using ACDS version 13.1 162 at 2016.08.22.07:15:55

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios is
	port (
		clk_clk                    : in    std_logic                     := '0';             --              clk.clk
		ddr_sdram_memory_mem_clk   : inout std_logic_vector(0 downto 0)  := (others => '0'); -- ddr_sdram_memory.mem_clk
		ddr_sdram_memory_mem_clk_n : inout std_logic_vector(0 downto 0)  := (others => '0'); --                 .mem_clk_n
		ddr_sdram_memory_mem_cs_n  : out   std_logic_vector(0 downto 0);                     --                 .mem_cs_n
		ddr_sdram_memory_mem_cke   : out   std_logic_vector(0 downto 0);                     --                 .mem_cke
		ddr_sdram_memory_mem_addr  : out   std_logic_vector(12 downto 0);                    --                 .mem_addr
		ddr_sdram_memory_mem_ba    : out   std_logic_vector(1 downto 0);                     --                 .mem_ba
		ddr_sdram_memory_mem_ras_n : out   std_logic;                                        --                 .mem_ras_n
		ddr_sdram_memory_mem_cas_n : out   std_logic;                                        --                 .mem_cas_n
		ddr_sdram_memory_mem_we_n  : out   std_logic;                                        --                 .mem_we_n
		ddr_sdram_memory_mem_dq    : inout std_logic_vector(15 downto 0) := (others => '0'); --                 .mem_dq
		ddr_sdram_memory_mem_dqs   : inout std_logic_vector(1 downto 0)  := (others => '0'); --                 .mem_dqs
		ddr_sdram_memory_mem_dm    : out   std_logic_vector(1 downto 0);                     --                 .mem_dm
		key_export                 : in    std_logic                     := '0';             --              key.export
		reset_reset_n              : in    std_logic                     := '0';             --            reset.reset_n
		led_export                 : out   std_logic                                         --              led.export
	);
end entity nios;

architecture rtl of nios is
	component nios_cpu is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(26 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component nios_cpu;

	component nios_onchip_ram is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component nios_onchip_ram;

	component nios_ddr_sdram is
		port (
			local_address     : in    std_logic_vector(22 downto 0) := (others => 'X'); -- address
			local_write_req   : in    std_logic                     := 'X';             -- write
			local_read_req    : in    std_logic                     := 'X';             -- read
			local_burstbegin  : in    std_logic                     := 'X';             -- beginbursttransfer
			local_ready       : out   std_logic;                                        -- waitrequest_n
			local_rdata       : out   std_logic_vector(31 downto 0);                    -- readdata
			local_rdata_valid : out   std_logic;                                        -- readdatavalid
			local_wdata       : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			local_be          : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			local_size        : in    std_logic                     := 'X';             -- burstcount
			local_refresh_ack : out   std_logic;                                        -- export
			local_init_done   : out   std_logic;                                        -- export
			reset_phy_clk_n   : out   std_logic;                                        -- export
			mem_clk           : inout std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_clk
			mem_clk_n         : inout std_logic_vector(0 downto 0)  := (others => 'X'); -- mem_clk_n
			mem_cs_n          : out   std_logic_vector(0 downto 0);                     -- mem_cs_n
			mem_cke           : out   std_logic_vector(0 downto 0);                     -- mem_cke
			mem_addr          : out   std_logic_vector(12 downto 0);                    -- mem_addr
			mem_ba            : out   std_logic_vector(1 downto 0);                     -- mem_ba
			mem_ras_n         : out   std_logic;                                        -- mem_ras_n
			mem_cas_n         : out   std_logic;                                        -- mem_cas_n
			mem_we_n          : out   std_logic;                                        -- mem_we_n
			mem_dq            : inout std_logic_vector(15 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs           : inout std_logic_vector(1 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dm            : out   std_logic_vector(1 downto 0);                     -- mem_dm
			pll_ref_clk       : in    std_logic                     := 'X';             -- clk
			soft_reset_n      : in    std_logic                     := 'X';             -- reset_n
			global_reset_n    : in    std_logic                     := 'X';             -- reset_n
			reset_request_n   : out   std_logic;                                        -- reset_n
			phy_clk           : out   std_logic;                                        -- clk
			aux_full_rate_clk : out   std_logic;                                        -- clk
			aux_half_rate_clk : out   std_logic                                         -- clk
		);
	end component nios_ddr_sdram;

	component nios_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios_jtag_uart;

	component nios_key is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component nios_key;

	component nios_led is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component nios_led;

	component nios_mm_interconnect_0 is
		port (
			ddr_sdram_sysclk_clk                                      : in  std_logic                     := 'X';             -- clk
			cpu_reset_n_reset_bridge_in_reset_reset                   : in  std_logic                     := 'X';             -- reset
			ddr_sdram_s1_translator_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                                   : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest                               : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable                                : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                                      : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                                  : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_write                                     : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess                               : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address                            : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest                        : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read                               : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata                           : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_jtag_debug_module_address                             : out std_logic_vector(8 downto 0);                     -- address
			cpu_jtag_debug_module_write                               : out std_logic;                                        -- write
			cpu_jtag_debug_module_read                                : out std_logic;                                        -- read
			cpu_jtag_debug_module_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_jtag_debug_module_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_jtag_debug_module_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_jtag_debug_module_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			cpu_jtag_debug_module_debugaccess                         : out std_logic;                                        -- debugaccess
			ddr_sdram_s1_address                                      : out std_logic_vector(22 downto 0);                    -- address
			ddr_sdram_s1_write                                        : out std_logic;                                        -- write
			ddr_sdram_s1_read                                         : out std_logic;                                        -- read
			ddr_sdram_s1_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ddr_sdram_s1_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			ddr_sdram_s1_beginbursttransfer                           : out std_logic;                                        -- beginbursttransfer
			ddr_sdram_s1_burstcount                                   : out std_logic_vector(0 downto 0);                     -- burstcount
			ddr_sdram_s1_byteenable                                   : out std_logic_vector(3 downto 0);                     -- byteenable
			ddr_sdram_s1_readdatavalid                                : in  std_logic                     := 'X';             -- readdatavalid
			ddr_sdram_s1_waitrequest                                  : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_address                       : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                         : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                          : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest                   : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                    : out std_logic;                                        -- chipselect
			key_s1_address                                            : out std_logic_vector(1 downto 0);                     -- address
			key_s1_write                                              : out std_logic;                                        -- write
			key_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			key_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			key_s1_chipselect                                         : out std_logic;                                        -- chipselect
			led_s1_address                                            : out std_logic_vector(1 downto 0);                     -- address
			led_s1_write                                              : out std_logic;                                        -- write
			led_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			led_s1_chipselect                                         : out std_logic;                                        -- chipselect
			onchip_ram_s1_address                                     : out std_logic_vector(12 downto 0);                    -- address
			onchip_ram_s1_write                                       : out std_logic;                                        -- write
			onchip_ram_s1_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_ram_s1_writedata                                   : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_ram_s1_byteenable                                  : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_ram_s1_chipselect                                  : out std_logic;                                        -- chipselect
			onchip_ram_s1_clken                                       : out std_logic                                         -- clken
		);
	end component nios_mm_interconnect_0;

	component nios_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios_irq_mapper;

	component nios_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios_rst_controller;

	component nios_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios_rst_controller_001;

	signal ddr_sdram_sysclk_clk                                          : std_logic;                     -- ddr_sdram:phy_clk -> [cpu:clk, irq_mapper:clk, jtag_uart:clk, key:clk, led:clk, mm_interconnect_0:ddr_sdram_sysclk_clk, onchip_ram:clk, rst_controller:clk]
	signal cpu_data_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_writedata                                     : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_data_master_address                                       : std_logic_vector(26 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_write                                         : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_read                                          : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_debugaccess                                   : std_logic;                     -- cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_byteenable                                    : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal ddr_sdram_s1_waitrequest                                      : std_logic;                     -- ddr_sdram:local_ready -> ddr_sdram_s1_waitrequest:in
	signal mm_interconnect_0_ddr_sdram_s1_burstcount                     : std_logic_vector(0 downto 0);  -- mm_interconnect_0:ddr_sdram_s1_burstcount -> ddr_sdram:local_size
	signal mm_interconnect_0_ddr_sdram_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:ddr_sdram_s1_writedata -> ddr_sdram:local_wdata
	signal mm_interconnect_0_ddr_sdram_s1_address                        : std_logic_vector(22 downto 0); -- mm_interconnect_0:ddr_sdram_s1_address -> ddr_sdram:local_address
	signal mm_interconnect_0_ddr_sdram_s1_write                          : std_logic;                     -- mm_interconnect_0:ddr_sdram_s1_write -> ddr_sdram:local_write_req
	signal mm_interconnect_0_ddr_sdram_s1_beginbursttransfer             : std_logic;                     -- mm_interconnect_0:ddr_sdram_s1_beginbursttransfer -> ddr_sdram:local_burstbegin
	signal mm_interconnect_0_ddr_sdram_s1_read                           : std_logic;                     -- mm_interconnect_0:ddr_sdram_s1_read -> ddr_sdram:local_read_req
	signal mm_interconnect_0_ddr_sdram_s1_readdata                       : std_logic_vector(31 downto 0); -- ddr_sdram:local_rdata -> mm_interconnect_0:ddr_sdram_s1_readdata
	signal mm_interconnect_0_ddr_sdram_s1_readdatavalid                  : std_logic;                     -- ddr_sdram:local_rdata_valid -> mm_interconnect_0:ddr_sdram_s1_readdatavalid
	signal mm_interconnect_0_ddr_sdram_s1_byteenable                     : std_logic_vector(3 downto 0);  -- mm_interconnect_0:ddr_sdram_s1_byteenable -> ddr_sdram:local_be
	signal mm_interconnect_0_cpu_jtag_debug_module_waitrequest           : std_logic;                     -- cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	signal mm_interconnect_0_cpu_jtag_debug_module_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	signal mm_interconnect_0_cpu_jtag_debug_module_address               : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	signal mm_interconnect_0_cpu_jtag_debug_module_write                 : std_logic;                     -- mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	signal mm_interconnect_0_cpu_jtag_debug_module_read                  : std_logic;                     -- mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	signal mm_interconnect_0_cpu_jtag_debug_module_readdata              : std_logic_vector(31 downto 0); -- cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	signal mm_interconnect_0_cpu_jtag_debug_module_debugaccess           : std_logic;                     -- mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	signal mm_interconnect_0_cpu_jtag_debug_module_byteenable            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	signal mm_interconnect_0_onchip_ram_s1_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	signal mm_interconnect_0_onchip_ram_s1_address                       : std_logic_vector(12 downto 0); -- mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	signal mm_interconnect_0_onchip_ram_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	signal mm_interconnect_0_onchip_ram_s1_clken                         : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	signal mm_interconnect_0_onchip_ram_s1_write                         : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	signal mm_interconnect_0_onchip_ram_s1_readdata                      : std_logic_vector(31 downto 0); -- onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	signal mm_interconnect_0_onchip_ram_s1_byteenable                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	signal mm_interconnect_0_led_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_s1_writedata -> led:writedata
	signal mm_interconnect_0_led_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_s1_address -> led:address
	signal mm_interconnect_0_led_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:led_s1_chipselect -> led:chipselect
	signal mm_interconnect_0_led_s1_write                                : std_logic;                     -- mm_interconnect_0:led_s1_write -> mm_interconnect_0_led_s1_write:in
	signal mm_interconnect_0_led_s1_readdata                             : std_logic_vector(31 downto 0); -- led:readdata -> mm_interconnect_0:led_s1_readdata
	signal mm_interconnect_0_key_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:key_s1_writedata -> key:writedata
	signal mm_interconnect_0_key_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:key_s1_address -> key:address
	signal mm_interconnect_0_key_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:key_s1_chipselect -> key:chipselect
	signal mm_interconnect_0_key_s1_write                                : std_logic;                     -- mm_interconnect_0:key_s1_write -> mm_interconnect_0_key_s1_write:in
	signal mm_interconnect_0_key_s1_readdata                             : std_logic_vector(31 downto 0); -- key:readdata -> mm_interconnect_0:key_s1_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal cpu_instruction_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                : std_logic_vector(26 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                   : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal cpu_instruction_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal ddr_sdram_reset_request_n_reset                               : std_logic;                     -- ddr_sdram:reset_request_n -> ddr_sdram_reset_request_n_reset:in
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- key:irq -> irq_mapper:receiver1_irq
	signal cpu_d_irq_irq                                                 : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:d_irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, onchip_ram:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                     -- rst_controller:reset_req -> [cpu:reset_req, onchip_ram:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                            : std_logic;                     -- rst_controller_001:reset_out -> rst_controller_001_reset_out_reset:in
	signal reset_reset_n_ports_inv                                       : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_ddr_sdram_s1_inv                            : std_logic;                     -- ddr_sdram_s1_waitrequest:inv -> mm_interconnect_0:ddr_sdram_s1_waitrequest
	signal mm_interconnect_0_led_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_led_s1_write:inv -> led:write_n
	signal mm_interconnect_0_key_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_key_s1_write:inv -> key:write_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal ddr_sdram_reset_request_n_reset_ports_inv                     : std_logic;                     -- ddr_sdram_reset_request_n_reset:inv -> mm_interconnect_0:ddr_sdram_s1_translator_reset_reset_bridge_in_reset_reset
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [cpu:reset_n, jtag_uart:rst_n, key:reset_n, led:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                  : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [ddr_sdram:global_reset_n, ddr_sdram:soft_reset_n]

begin

	cpu : component nios_cpu
		port map (
			clk                                   => ddr_sdram_sysclk_clk,                                --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,            --                   reset_n.reset_n
			reset_req                             => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                             => cpu_data_master_address,                             --               data_master.address
			d_byteenable                          => cpu_data_master_byteenable,                          --                          .byteenable
			d_read                                => cpu_data_master_read,                                --                          .read
			d_readdata                            => cpu_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => cpu_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => cpu_data_master_write,                               --                          .write
			d_writedata                           => cpu_data_master_writedata,                           --                          .writedata
			jtag_debug_module_debugaccess_to_roms => cpu_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => cpu_instruction_master_address,                      --        instruction_master.address
			i_read                                => cpu_instruction_master_read,                         --                          .read
			i_readdata                            => cpu_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => cpu_instruction_master_waitrequest,                  --                          .waitrequest
			d_irq                                 => cpu_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => open,                                                --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_cpu_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_cpu_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_cpu_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_cpu_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_0_cpu_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_cpu_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_cpu_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_0_cpu_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open                                                 -- custom_instruction_master.readra
		);

	onchip_ram : component nios_onchip_ram
		port map (
			clk        => ddr_sdram_sysclk_clk,                       --   clk1.clk
			address    => mm_interconnect_0_onchip_ram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_ram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_ram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_ram_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_ram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_ram_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_ram_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,             -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req          --       .reset_req
		);

	ddr_sdram : component nios_ddr_sdram
		port map (
			local_address     => mm_interconnect_0_ddr_sdram_s1_address,            --                  s1.address
			local_write_req   => mm_interconnect_0_ddr_sdram_s1_write,              --                    .write
			local_read_req    => mm_interconnect_0_ddr_sdram_s1_read,               --                    .read
			local_burstbegin  => mm_interconnect_0_ddr_sdram_s1_beginbursttransfer, --                    .beginbursttransfer
			local_ready       => ddr_sdram_s1_waitrequest,                          --                    .waitrequest_n
			local_rdata       => mm_interconnect_0_ddr_sdram_s1_readdata,           --                    .readdata
			local_rdata_valid => mm_interconnect_0_ddr_sdram_s1_readdatavalid,      --                    .readdatavalid
			local_wdata       => mm_interconnect_0_ddr_sdram_s1_writedata,          --                    .writedata
			local_be          => mm_interconnect_0_ddr_sdram_s1_byteenable,         --                    .byteenable
			local_size        => mm_interconnect_0_ddr_sdram_s1_burstcount(0),      --                    .burstcount
			local_refresh_ack => open,                                              -- external_connection.export
			local_init_done   => open,                                              --                    .export
			reset_phy_clk_n   => open,                                              --                    .export
			mem_clk           => ddr_sdram_memory_mem_clk,                          --              memory.mem_clk
			mem_clk_n         => ddr_sdram_memory_mem_clk_n,                        --                    .mem_clk_n
			mem_cs_n          => ddr_sdram_memory_mem_cs_n,                         --                    .mem_cs_n
			mem_cke           => ddr_sdram_memory_mem_cke,                          --                    .mem_cke
			mem_addr          => ddr_sdram_memory_mem_addr,                         --                    .mem_addr
			mem_ba            => ddr_sdram_memory_mem_ba,                           --                    .mem_ba
			mem_ras_n         => ddr_sdram_memory_mem_ras_n,                        --                    .mem_ras_n
			mem_cas_n         => ddr_sdram_memory_mem_cas_n,                        --                    .mem_cas_n
			mem_we_n          => ddr_sdram_memory_mem_we_n,                         --                    .mem_we_n
			mem_dq            => ddr_sdram_memory_mem_dq,                           --                    .mem_dq
			mem_dqs           => ddr_sdram_memory_mem_dqs,                          --                    .mem_dqs
			mem_dm            => ddr_sdram_memory_mem_dm,                           --                    .mem_dm
			pll_ref_clk       => clk_clk,                                           --              refclk.clk
			soft_reset_n      => rst_controller_001_reset_out_reset_ports_inv,      --        soft_reset_n.reset_n
			global_reset_n    => rst_controller_001_reset_out_reset_ports_inv,      --      global_reset_n.reset_n
			reset_request_n   => ddr_sdram_reset_request_n_reset,                   --     reset_request_n.reset_n
			phy_clk           => ddr_sdram_sysclk_clk,                              --              sysclk.clk
			aux_full_rate_clk => open,                                              --             auxfull.clk
			aux_half_rate_clk => open                                               --             auxhalf.clk
		);

	jtag_uart : component nios_jtag_uart
		port map (
			clk            => ddr_sdram_sysclk_clk,                                          --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	key : component nios_key
		port map (
			clk        => ddr_sdram_sysclk_clk,                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_key_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_key_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_key_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_key_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_key_s1_readdata,        --                    .readdata
			in_port    => key_export,                               -- external_connection.export
			irq        => irq_mapper_receiver1_irq                  --                 irq.irq
		);

	led : component nios_led
		port map (
			clk        => ddr_sdram_sysclk_clk,                     --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_led_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_s1_readdata,        --                    .readdata
			out_port   => led_export                                -- external_connection.export
		);

	mm_interconnect_0 : component nios_mm_interconnect_0
		port map (
			ddr_sdram_sysclk_clk                                      => ddr_sdram_sysclk_clk,                                      --                                    ddr_sdram_sysclk.clk
			cpu_reset_n_reset_bridge_in_reset_reset                   => rst_controller_reset_out_reset,                            --                   cpu_reset_n_reset_bridge_in_reset.reset
			ddr_sdram_s1_translator_reset_reset_bridge_in_reset_reset => ddr_sdram_reset_request_n_reset_ports_inv,                 -- ddr_sdram_s1_translator_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                                   => cpu_data_master_address,                                   --                                     cpu_data_master.address
			cpu_data_master_waitrequest                               => cpu_data_master_waitrequest,                               --                                                    .waitrequest
			cpu_data_master_byteenable                                => cpu_data_master_byteenable,                                --                                                    .byteenable
			cpu_data_master_read                                      => cpu_data_master_read,                                      --                                                    .read
			cpu_data_master_readdata                                  => cpu_data_master_readdata,                                  --                                                    .readdata
			cpu_data_master_write                                     => cpu_data_master_write,                                     --                                                    .write
			cpu_data_master_writedata                                 => cpu_data_master_writedata,                                 --                                                    .writedata
			cpu_data_master_debugaccess                               => cpu_data_master_debugaccess,                               --                                                    .debugaccess
			cpu_instruction_master_address                            => cpu_instruction_master_address,                            --                              cpu_instruction_master.address
			cpu_instruction_master_waitrequest                        => cpu_instruction_master_waitrequest,                        --                                                    .waitrequest
			cpu_instruction_master_read                               => cpu_instruction_master_read,                               --                                                    .read
			cpu_instruction_master_readdata                           => cpu_instruction_master_readdata,                           --                                                    .readdata
			cpu_jtag_debug_module_address                             => mm_interconnect_0_cpu_jtag_debug_module_address,           --                               cpu_jtag_debug_module.address
			cpu_jtag_debug_module_write                               => mm_interconnect_0_cpu_jtag_debug_module_write,             --                                                    .write
			cpu_jtag_debug_module_read                                => mm_interconnect_0_cpu_jtag_debug_module_read,              --                                                    .read
			cpu_jtag_debug_module_readdata                            => mm_interconnect_0_cpu_jtag_debug_module_readdata,          --                                                    .readdata
			cpu_jtag_debug_module_writedata                           => mm_interconnect_0_cpu_jtag_debug_module_writedata,         --                                                    .writedata
			cpu_jtag_debug_module_byteenable                          => mm_interconnect_0_cpu_jtag_debug_module_byteenable,        --                                                    .byteenable
			cpu_jtag_debug_module_waitrequest                         => mm_interconnect_0_cpu_jtag_debug_module_waitrequest,       --                                                    .waitrequest
			cpu_jtag_debug_module_debugaccess                         => mm_interconnect_0_cpu_jtag_debug_module_debugaccess,       --                                                    .debugaccess
			ddr_sdram_s1_address                                      => mm_interconnect_0_ddr_sdram_s1_address,                    --                                        ddr_sdram_s1.address
			ddr_sdram_s1_write                                        => mm_interconnect_0_ddr_sdram_s1_write,                      --                                                    .write
			ddr_sdram_s1_read                                         => mm_interconnect_0_ddr_sdram_s1_read,                       --                                                    .read
			ddr_sdram_s1_readdata                                     => mm_interconnect_0_ddr_sdram_s1_readdata,                   --                                                    .readdata
			ddr_sdram_s1_writedata                                    => mm_interconnect_0_ddr_sdram_s1_writedata,                  --                                                    .writedata
			ddr_sdram_s1_beginbursttransfer                           => mm_interconnect_0_ddr_sdram_s1_beginbursttransfer,         --                                                    .beginbursttransfer
			ddr_sdram_s1_burstcount                                   => mm_interconnect_0_ddr_sdram_s1_burstcount,                 --                                                    .burstcount
			ddr_sdram_s1_byteenable                                   => mm_interconnect_0_ddr_sdram_s1_byteenable,                 --                                                    .byteenable
			ddr_sdram_s1_readdatavalid                                => mm_interconnect_0_ddr_sdram_s1_readdatavalid,              --                                                    .readdatavalid
			ddr_sdram_s1_waitrequest                                  => mm_interconnect_0_ddr_sdram_s1_inv,                        --                                                    .waitrequest
			jtag_uart_avalon_jtag_slave_address                       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --                         jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                         => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                                    .write
			jtag_uart_avalon_jtag_slave_read                          => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                                    .read
			jtag_uart_avalon_jtag_slave_readdata                      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                                    .readdata
			jtag_uart_avalon_jtag_slave_writedata                     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                                    .writedata
			jtag_uart_avalon_jtag_slave_waitrequest                   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                                    .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                                    .chipselect
			key_s1_address                                            => mm_interconnect_0_key_s1_address,                          --                                              key_s1.address
			key_s1_write                                              => mm_interconnect_0_key_s1_write,                            --                                                    .write
			key_s1_readdata                                           => mm_interconnect_0_key_s1_readdata,                         --                                                    .readdata
			key_s1_writedata                                          => mm_interconnect_0_key_s1_writedata,                        --                                                    .writedata
			key_s1_chipselect                                         => mm_interconnect_0_key_s1_chipselect,                       --                                                    .chipselect
			led_s1_address                                            => mm_interconnect_0_led_s1_address,                          --                                              led_s1.address
			led_s1_write                                              => mm_interconnect_0_led_s1_write,                            --                                                    .write
			led_s1_readdata                                           => mm_interconnect_0_led_s1_readdata,                         --                                                    .readdata
			led_s1_writedata                                          => mm_interconnect_0_led_s1_writedata,                        --                                                    .writedata
			led_s1_chipselect                                         => mm_interconnect_0_led_s1_chipselect,                       --                                                    .chipselect
			onchip_ram_s1_address                                     => mm_interconnect_0_onchip_ram_s1_address,                   --                                       onchip_ram_s1.address
			onchip_ram_s1_write                                       => mm_interconnect_0_onchip_ram_s1_write,                     --                                                    .write
			onchip_ram_s1_readdata                                    => mm_interconnect_0_onchip_ram_s1_readdata,                  --                                                    .readdata
			onchip_ram_s1_writedata                                   => mm_interconnect_0_onchip_ram_s1_writedata,                 --                                                    .writedata
			onchip_ram_s1_byteenable                                  => mm_interconnect_0_onchip_ram_s1_byteenable,                --                                                    .byteenable
			onchip_ram_s1_chipselect                                  => mm_interconnect_0_onchip_ram_s1_chipselect,                --                                                    .chipselect
			onchip_ram_s1_clken                                       => mm_interconnect_0_onchip_ram_s1_clken                      --                                                    .clken
		);

	irq_mapper : component nios_irq_mapper
		port map (
			clk           => ddr_sdram_sysclk_clk,           --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => cpu_d_irq_irq                   --    sender.irq
		);

	rst_controller : component nios_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => ddr_sdram_sysclk_clk,               --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component nios_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_ddr_sdram_s1_inv <= not ddr_sdram_s1_waitrequest;

	mm_interconnect_0_led_s1_write_ports_inv <= not mm_interconnect_0_led_s1_write;

	mm_interconnect_0_key_s1_write_ports_inv <= not mm_interconnect_0_key_s1_write;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	ddr_sdram_reset_request_n_reset_ports_inv <= not ddr_sdram_reset_request_n_reset;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of nios
