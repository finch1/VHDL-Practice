��/  ��^k*��A��D@7�քW�g̝�G�^�T�|�IVϪ�y�p;�5��p:#�oj#�_�����H�+k��'O 5aj�[��l��Åéh�?��dDH�ݻy�RZӢXbf�p���xmt�[+hH�1y�
o��C��%d]���Tz����q���x��Q%MM��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ��W�Q��L�Uт�X"��ؖ��1�O[�B���:��B�X]U%�n�g��5����͉�׃PuO�]��p�>6BD�d����MNM�è�%���*Mw��s?v5��P���]�]�$������[�>.��a��B,�g��Lð�p���f[����R��ix�b��B�?�o�r�hV��L^GR��zҀ�C揻r�K�\�>����q)u͞����m&�(��G�FY=�����ߝ�@�b`�*�{`�3�n ��K�31���G�g�r�1�Gvd{�t+C�X�J��\P뙏�lBO��9�����s`���e��q�h��c�?*y˨���HI��h�>��R?e�YExgU!�Z�C�>!�S����R�Vȼ��K�V�=<��A��%��[8ʔe���k��*H��ej�h���X�R�n�DY�%�zp]\�:]7����D5��K�2�nWl���zf�����*�9�K�� �Jv����`�A8,�ڂN"�E�� q��<�ɭ��"a�Wx�/�~��h��V��<Մ&֊*���/ w����c�
����p�C���37~�DvQ��vh��(Y,1M:b��8��t(�E�C1K��a�����~��
�]¤���#������K�8�ǐѲ�t���n�du��ZP�ZB���UgP>���g�Y�x��Oa,�������u� >6��)Ѝ ��B0�]���#(ֆ��x����y�:.!߃8���RJ~1�w�8e�LO�!�dAKa�y3����hA���şlY�v/4T���1��wש��R
ߴs׌���t� ��;��]��LfÄ'�S����6�r�=�F�>��tW���Z��;$����a���-k��V7T2��!g��3����W���ll�g3�� n���:����Iς�~�p_��X�ƨ�3Bt����rO��3/6|�	 ��hl�˰�U�a{�]+v�!:!�Ńˑ?C�c4�	T���ef�o�;�ؿ��Sr�69~�˲��Hwe��"dp�ș��D:�I�2i1�I�,�2JQy���9�k\��Cl�P1�H��F"k����Gh��e��)�)B�CB>
0�Kߦ�s}�1-��uy��pE�ۑ��"�8�ϔ|R#츭_�x�'��B��jP��Y�I���ᮀ�#������ CN�!}�N2��g�3�v?Q�b�U����g��IH����)o�� �l�Y�p��ø�7��S��Jls�V�u:��1}6 �Q$�}�ٱ�0��Y�X��H��hP�C~QP�CH<�ǗW��jȖ�횇���h�IRbn3��]��uW��3�OP ��ayJI�Q�-F���nŚ2�=1Z%����j��'O'���I�|F4�*����H�̑O_�{� �gu�A
�W2
(�tT_T5�-���z�ПZ΍��� �Yy�mt���2�!*����7Bv$�$$�c/^u����4M�rT�O*�!�Ƣ#�k�A��y��q�g�{�P���n�f0B�eQ.�*���	]��p��e�O&w�r��=K����:�CzI�J�ąy�������P��(��۔)���Wt��ȗ|B�5˝vz�Q�L���gԿ�zS(8]O����&�f;Ѓ$���_�W-�n��ov:7pu9u#/�	���h�{O�D��B���q|���'�����ł^0�)p��'�n���ce�t��]u]�[�������,g���Ⱦ��(�e�:hm�E�J�۬�/�<�O~�4s<�,���(l K�~V.��M���EG��SVLz�Ze���4�m<��4惔�B�� �b������޶���;��玶I�Ы�
,���ە:�c�TC`rL�"�I�Ŋ�X��/=��(i�l��4��(}���_�Q�l��諚��#e�7�s�Ћ �^٨�v�Ǵf�������K��i:��x >�pr�dr�ɑ��0hК�b�1zs�P�[� >�^��\~;�����m������7^�u;|���_���^R�-G�O]�C��!��]D-6�
NSؒ
�Ulʭ�U��D�*�i$�IK�vg��U]��G���?A���������r����P��-��)�=�dD]"�t=jZ�m �PN�p�u-3��H���x�E������]Z.-b��r�r��i��s�x.�� ���b��(@�ݷ��b��c��mO��p)�(9��S�M`N�u�ZL�Ӛ�,9�?3eB��J+C���'*\t�����V���'��?E�]�`S>��n\{˴�!ĽY2��y�����S���W�w��|M�`Ź�HZM�D5�^����o�v��KрD��>������.f}y�.�u�c]����R���C|�h�۹���xvk�f��� �k�b�J�m�{�������N1�Kw�*�vp��X�s�0�h�}�l�	��)���='�C8�|�s@>�P��@k:*��Km��o�2IQ$sV��l�k�Q;�
��T�M�K�_g�}߉4�I����(���i�أ!��49+A������Ý���+&H�0ar5��~��Jڒ�E�"��ct�6���m�a��0��?�.�����*"��|�$�h���3�j��؁���������6������Ǣ��	��	�uѯ{��~�TQ�k��6��M*���ꮒ?��Ƹ��ϯT�Z��4�S�h��	�f
�afi���?xQ�!�J\��>-[��T*��e�5x}Yv>#}�ѥ1�!������E/M��� � j��+�^d�]f�y*�=P�J�A�2Y�`��c�|��ש2�6x�"��j����	�ݺT�Q�Zs[�/ԿER3j>�������� ��硞�;��*�,g*�#�F�ƝOr�T8��&�P{�?���ca��KD�/?��l�*��S�A���sZN -2qX��V(���������B1.�v+�Ub�o�˲&����!1�m�;�߈�h���z���<�j$�[�x�F-(��GMC�T�W3E�����\s��&5�h>i[` GTU��>��h�U��qɎ�Ƅ�?�Q�����*�8!>�n�-$�; �m�O��?�7�d(��Y�}�"��Og%�-]b���^��!�?*R2a�"yl���7� ꪆWi�u�ӄ�G�/|(�HF�#����6i#���J�>���)#��Fj�$�v�B�/\E�3���d����ѓU�Q�B�� VB|�5���)�s%L�`U�'	���S�(��p��$��K���2�+�@�v'Cu��?W��R��:i��\"��7�� u%[��d�q^��R
��gz�E�e�_Q���8L���<�K?����Шل�\0y�f�'k{�"=����<�.5X���:(g���W#�K"�{זG��l�v�����HF�p�է҈5vJ1�3N��Xm�U�NN!�|�`������t�'��:K�5���0U���;�cp&xܠ���PKճ/t���Ma�\������]p���t�j�3�B��^�O�O���jn�R}߈�\ķ���:�w 𿜦��K4bٱ�7O����޵8��Sx�>l�����f�8��E0������`�R��Ȍo�>T�*l�8���U�s����t캗,��i++�h��ͽr���"� ������b<Kڡ�u������#�쫶(�_�34��D�R�Svx���<<f�B��qW����d�$���4(�NX�LTt��*�/�b��qd�G�hm�fy���]���������l�sH�6��/4��$�w;��䅆�x������y��f����!A-�����=Jե���#����ɜ���Z�AQտ�9\:�������8 >��n�ڵ�x
1�j~�{`�c=ܭ<�����o�5c����/My��2��m]�Yh�6�MN�����X�-'�$hL����̧��G]eO�o��S"�c����0�A�H.-���ہHُ���,P�,C3��U�ZzH+�s �F�}4�x�D�V����p(�3)��H{�i�9D��������$��{�ZQ����%R�����_ʨ�=I�h!\{Y�^�j!�%�$0�����hb���d�E��
d#Ѯ0���>�ݎܐ<N�����J��-��(��;Y��O}[��lТ��>�h�b�>_$���1�V�����~���O��t��~s����1d:�p����نb�buE��/	��s��r���;�3D���Wq\Hh��z��I�*���J�5�z3��͢�@��	���'f��{�ͬd*Ѡ�=K&_�_���'�K��ڏ��RP#�>���%F=�~.��a����Rb����K�S�;��%2(�Y��l;����l���|������DT�p��ul�貶��L^���E溙��n�q��#$�Ȥ����XZs��^C���'���!�H/B�S�n��U^➴���e����"��VN��5�����D����������b��R�ĆK�y]a��cY�>��TÜ�;��@ ��	�=.@x��Ԃ��Ð��Ӹ|��n�"%���ņ��������;�	���e�ژ��qټ��={�9�)_�2������{_.�z����@�?���O�����Bw��r��5̗�Ɖ����ٙ)�x� �apy',J}sS�l,+�cR�[/��_�8?sQځSUa���zAߞ�g];��G�!֡�`z�(:�gyr`�����fM�ej��H��J�%L�+E���:7r3F)������/�"�����YL N}(���O�qM���U�ϢQ�ޓ�4�`,��`�P���`m�wQ�)[燂�Ջ��1�F�qcy��S�㥇�=C�f��@�O���<���R�B�J�gf!��h�6�G��1�1�h��pojd�:ypb��+���9[��gJ�k"�1��*G�t�-�N�c�N�
�9�ͩ<Nh-�5�PT2f�^��^1�3�ڷ�q����O'�g�=N����	�f���Z�����t�ǘ���~��4/�s]��=�������kZ����3�(��|P*�%����#�;�ż��X2� ���Vc�e��y��rO���������$�n!�'BHI���S�`�-\�
����/����	��4�@���u2�O��m2�9�ƍ�u�Ъ��ӭ�M�]��>�i�N�܄��Z�~��0�Q_��R�omV�@h�_]��O�e���$�D��#��1I���8�9��f�<��ݔ4Fм���ѻ-��!����{��S�b��	X�#��q��O��w��(��8U�4A����%�W��]��v��-.�Z�'��}�p��H�r�41S
|�F������`Q��}E�����a�g�ė`s����I�O����Žc`bM=�sc�3��-Gȩlg�%�a���*^�V�i��1����^���}����������tQ��J�mc��|�}ko��E�e�#���s��ݼ�G���yh1b5P��M8��>T�v�|j����]�/n\d4�Y5��2�~�i��>X�:�M�j3����W�M�T���Wf6X��.�^��(�MGDWl�\���#�"i��lk"%-Z[J����U���-T��g��~;�$AV���?��Y 0� /�T$m�t&�/��f;2�t3�ܡ���z&�����W�@c@^.�buF����+XD����bn���[�r`�5x�n�q���8�%I�+�$��T_�\l���ڬvL��+���Y�E�����/r��>�ւ�1n������ظ�%~U��W�u�'�RC�7�"���5�喣�ğ�=����K�5v�7��\uf+��t G;���o���`��x��X�)����5oU6��'��D�s�>��
]��&�P�1)Ь�b7�q�[:՜����U�Ɗ�jf���a��{��,�z7������<JSC�>YP�ݜ3 ��@�6H	�i�T�������T􋣆�Al:cޒj���C�N���H���
��>3���^��'n��J�Kl�x<N]� ���������H*$���Z�B�����ԃ����"��?��F��4��c�B�h+����	���a9���6TuG{xV�6�[R�����)����[u�O��47р��.�9h$�k���=���N��#1�7�h@pzf��h��N�	y9 R,���l3��ˎٛ���ʢ²�q�.�9�7۪�7���z�i��4e �9�|h������ �u��R�Hd݌��1
S��qa�6�iN���?��]�ê�O��%��,�^��D;��8�����y]�Y+%;��N��O� 5�]�\�f�Q�2:l�K�·k�I6&��Gid2f��'떓�LK��?0�3Y���g��� �#��ON�׮s/��$�$;����:��)��1I�~F�+F���5��Ụ���/��?AP0���J�����y���<ح���Z��v�z���p@�-yꛥ���$�� 57$ S���#Wm��VG���t������얼qR���&���.!�t5��:?�! �M�}�>���=�>��R�	Ϣ/��ltG�qզ��~<X)��0;��HRެ��W�ź���0$-�0d����T~�@�ⵊmb�f.n�n:61P�Hs�8fo�a����Uj�����c��g��?��
f$j&T�4�˿�[!Q�ǚ��~sԨsߐHO^#��bM%�H�S����=�f���K�џDwOE���
����W�\]a�.�3 ����4���pY�R|�fs"��7L����/Ŝ?��I� Ϻ0��b{�[I�JК��KFiI	S��%�E�`��n�$3M�?y#.���c �I����reK��7G��or�
�^�1-gB��;E�U��4X� i�i0��c���)v�C��� ��J�1���m����w�%���p�Dy�'pN&'�2��@b�Ym�OӨN�=�fg-�'Nӊ�r�ɱ���nAJ.-�,���`�lཥ_l��|�ӻW*:���B�l���K�,�6����-��P-����n��Y��C�R�)���i=U��v�|����3 ��=_6�c/3Ҿ��x޿�W v�F����k��`$�s��T����t���AlH���s���k�N;�*C�f��|Y���P�9��`��� ����-�u��%Y԰F���x��Qa`Γ���U�ǿ*�$�޶>�$.T!!Ԇ_�֮�]]�ٲ�Udb����V��o��W�ׇ-k�d����E�z�ŋy:��
�i��(������������>Lo�	�}In$7(H�M��kU�
"���ԩ�$�@�dZbF��8S�q\�E������9D��3OJo_��b#������Rj	Nc��A���jTR�#q��|N�?+�s�e\Pi���(��h�Fw����Y@]��z�"�������k�õ���M�o��#n/�if�r(�=b�^j|D]��l?�!�}]��S$P����	�����R�����!��)�<�B�X��� ;�Ct���Œ,T0��x0e�ߕk ' 9^��+	z�yrr���~퉚T�rF�5��u��&j����'���*�	�g�_n�}U�d2����Ui���-��`T��o:�`F��bg���� @���o����q:�4���i��0��ǅ^�0��TzU���焒��Բ$�	�n����U�AS߻:_��8��"��>e�Mm^��JЪ���Z�p"���#KHb�?|��B?���&����.f��@]�?��!��Z�_�:��No[j�|�k�	 ���W/n}#6���h���,
�����m�Bg�����`�r�(ݴ�,����Lt<Xaֿ�)���4G[=2�ِ�z��)X�	��s�V�1ȦVY�yျ� 9����=�s<������f����d4���6���k�R�#�G0D���ܛ�[��v�4Tj�w_��Tc�Ijz[ɴM��<*�o'C֎�1�kC�fF�YB�oJ$�x��䰙�?�J>�4��3�1�"� uG�+�oxɥ�	�fx�Άs�#�5�e������]i�,&R��+:<�.�\�3:S���\����@���:�Ϛu�m�n��]Z����[B��c����H����z�f�5��V� h7;�1E�7�7����#�d7H�U�aCy�N���%�t×4��&r�?��#���X�X̡��8��?�>��vW֚�WUr�ʾɀ[��ŝ���RG/�}f� �b�s�ն͹���ؚ���B�H!~d��*ZH1�I{�Ak���0�7C���n��(1�-�Ȧj�o}�%w[��H"I�~Xw��s��d��GS�:"W1;��p^����&�A�x"6�V�U�t"�2,�s����m�\���Y�����k���4r�����M?/,k�2��i�Y)�m
���_���W�]YW��&��Ʀډ,��٫�k��9��D����η�|3Zԫ�E�39�U���\�ڗ7p�Gm��O9\.��.�:M�oת(m�&e{M�� ���f�IPK�O��t��V>x���)oCM�tz�{feyj&��q<��>�D�E[�l}�`�b��>�	�=6=M�D�W��u"�O[�{E�.h�ٯΠ�B`��?abK��<���u���؊@(�e+AH��&�|�*Z�8����z��\�����G��BahL�0wV���4Y�g2X�.d@�*��f��;���_��C�4�����kY�I���}�o4AV�3��F�ʻ�c�{�%q��~�<���4v��MǍ��y&�h��Qlr¤�=e�
����N��z��: ȡ�y�V�����8�i4�@�w<����?�i�j�?��VI3j���X�U��~����h8A�4kZD~�����nqt��c�
^�����p.�Zc����Gv��s]����ю�Yp�#�9%��Y�^d���iY��6�om-� ��o/�|8�h�/�
d�G�f\����撜)ڋ!�?���# 乄��[B�e�p!�1�U.
�6@����p�T#M��#K��������c���T�Ɨ��I��q%bsS�o£�(�z�薪������Jc.�e��DX�0�֬F���&۾3#��S!�ʯa��	v�9l?�c�O��
�1��������v+EGhc�=>�ٯC']�0h�$[V��Xi�A��qL���Ȅ�Uw�������M��)W.��ߙ ��}�S��ɍe"�c���Y���x] ��$�H�"�ɲ�I��[��3"	�����OV�*�}�|��fO!xD��<T(��O�{�Kj|��4,�� �'��k�٩�*��Pgr� T,��P���Є�P�T�`o�}�bI]������]T����(�8�8�����OBOdS-���1��c�C�vG�]IT�yN.���&��wB�N�(�IM�ǩm}�@�����$;g^b4=�y�:O��H�@������wC��)�=ã�6�)�C'cG��{�Qzb�E�/��FŖK�Y��)��R '�0�g|���Z6u�����ݎ�%�R��ð�P��3~�s�M�<i�<�O�YVQO8FG�H�?h�9��"��jO�\W=,��b4�� ;7��!
%�Cg�C+�r��x4���=�}��X�k��Pg���))y/�=���TXd)�E#`���%w���5���8�G(l>�vE��X�sG�?�u�!1��\�7������'3�<"˹��ř��펥j����w��-�`�cK� ��SyQ]�w�a\7�ӑ$��<
Y�~�g�|C��Y�NZ���TU�;h0{Ga�m3c$�\���}fX��dep`�1��r�e3������
�~y�qΈ�
�5� ��(�����^�b�������́��Ω�Ίp�X��},�
�	+.Ԭ/��W[�a�d���ʰ�*�5�T�R�3�ʂ��	
 �8�c��,T`W�;�9���W0K�,�������t.9�.i&��ў �o��������7�u`Y�\�pl#g)�]d��d�?����T��/�Ya��M�'і�������+�ɔ���xYڛ��`�Ky�I�'��bǡ�F/��/#:����o#<AwK�3	j�ɠ��(�p�n��Ǻ7$U$��x5��^���س�(F�,���⁕'���tjV��[DH�W���m�U�)o"6άl���j]��Gn��i�f�1׫��vz�4G���/+��{�2� �T>���}ל�1�Ru8��{���q��bٵ��W1Uk,�`��#�CA��|]�㯏}��>��rY���.��J�ϣ�r��ѫ6ׄ���i�Ԛ�����l��{���yTN�Xg�깮)��a$w�XZ���F��E\��Lp��:��* Q6N��[b���1;�*�"��j���%;+d�8��֛�*�Z c\�do����k������N���kr�x(f1(N�44�H�8+��X
*���++f�*��`��2�,�B�]z=�ܷ��\��4>Y��n�S�"KtOt&L��g5��b��j���ٱG��:���Tm0�-�%�4;������>�Y՟'+r���X� �ͮ;���A�@�$b����mbH�%|z����W�az�3H����g�8���������߇�ଫ+��;V��k�� �~z�YFD���ŋ�Hֵb��(�9SQx}�r'c�݀��䛪�br#��.�]���חܙ+�+�w��vθ<��W�C��z���--��UX����m��W��
k�Kl\SP������^���jm��7X71+���^\OWp��N��J�N6����q��� �uF�|X�{���YX�����V{"aD������-���h�Ə+� +n�Qkޮ�?E��0��"n��3���-1�㐶黍�MsdExzH��P~F�� 2<u��A�<zM���X����NhYR�ӷ�����>oaGP�"�s%�A��B��`n�4���=:�ww}R��]�����9(����\W{P���z�Z3��ݫ�{��Z��J]��9��8����W�Y�iE<?���T;�HPjz�0�z)�mGf�<�(Ýɠ��W�a؇����'���gM6[�g���:ۆ���_TJ!�Pvb"��O-����K�Bvl�\��m[̂Iz>�JD+ �������˥��D���������O��H�+/X<V��@����|�N���>���d���Ȭn���j�v�@U[<x?����4FT�� �k�bz�ԩ?ɳ�>.�j���v�:�k���$��r*�0����_�^T�]}�} ��a�[�0���CA=�2�i����̄�Ns�n�s�;Ku`�k����|��*1ّ���{#��-�L&�3p�k��eS]�i̬Y&�#)��O�ROr����w�b���8�k���01s疥��5������1fm{�o��}_N�"�t�m����g������;�� ���F�eX�����"z%O�����-����S0��~RW'����,ߤJ�s�vp]J'��0Չ���/�T�����

�<�U7�/�u�Ekj��>��.$���DVy_�ɔ�7�7�L⪠L�^A��=1�ȃn�&�l�4�.����j�������(��8��b#p)~4��22��'�ob�Δ��b&�iA��2!�V�^*��W��F1��6�>�~ޏ�s+��ƪ�γ�+A:�I
X�n���K+�Z��?�9���7��4?��Ǆ� �n�n��������p��%���ɦ��ٟ�W�w���eڿU�+��K~��o��i.(3VkT�#)J5��_-�CZ�������Z�1.C�SR����N�@=m3�?[J���7~L+��m����I�ACܦ��ؕoP����� ���
�?[}?1V��&=� ���
�6�BK�c'j��K݊n����H�����oH�C����n�(���I"j��\a�0�,�,.02�K���m��W������l'F�
�nQ�Ft-�1p6x
T�:���\���r��W~�m���4�����l��ޙi�qz�8%~>��8ɲ��4�6�ր��#ʶ�ں͜*�Hi���b�[b��K��i�B��~�Ϗ7d:<`D���J�B���󏈗�.aܘe]����ٵ��S���O�v>
�Qv�=u�����I�����	�Bw�����tc�$Y
�G��iP�<��v'��i
���=�o� �N��o�Wڂ�z*o ɕ�2�\lF,�xP �h�d�E�$���63��m����zB{�\ˋ�W�Œ~0[�q�ձ�W)�Oh0�s�2��$0�阥�Ҟ�W打E��=����ϥn���Q�vc�:��q�.���[Mۂ��g�]d��n�W!�KѿV���$�ϊ����e�+��3���������l]s��S���X*�[���U�~Ŵ��ț��4�jRD�~���w��W����ͩ0���-��	-��c��a�Qc�-(ψa[s_kuX��@ݷ],�m�B���2i't;'��LX�^��b'c�=1}���ˋ?�0�Qw��Bl+W�F�_�@x��3bP��#�N��>�M�Фw�=O�6����c�l�^��?�ɩ��$?"m�U�&R�w�tU0���w-G� 6�����6^�G����@dE�D�Q�B\�_��#��
=��4[���>�V�h�<������\�^co�AU����0����NR�)p~{�J(&��՜��oz0�CL����>,��NF? ���Q3"����4�09�� K!}]���@b��xdna�s��x$i�/�L���w�k��Q{��3]��/˲�h�C�lE�z	O~�G�X���+U%�(7�p�n���?����2(�̨;n�#�# ��h�v�]��h0���'cE�p�n7��Уv��+Q��-;�,vǥ��7�׹���p�_o�� �EVq���vP��)�i�̏&Y�\���d����˹������a�����Z՝�ׇ2J9���j�C{E�����������ۧz�ʞi#�ֻ����ÀN�J�����u
J�zm��Q3�[����d7��w�9(��h�)��֨|�ᯃ'Hn�,�K���j!�ԓ�^ҝC�7	t�[��*�yC�K�MY�'E����OLM�� ʙ��"!`�0#y1��ր|�ݸtd��2��VH�LG`J5c��/�p��g[Go���j���=L�9AN�����Ih�V+_���x���H�o�_����0�uB��
������m�M�We�3<]�6G�j�u���&.Py�'��#, ��c�ImZ6�#��"��Ȅ�4����E�l�"����.��(M>6�xi�M拏�^���}�6O���|8g�v�Q��o�u�6},Jj8���WƲT��w!����0��^��>��K�卝�Ζ���si˅m�o6Tw⃝ohj�p�apk�J����4��j�����������%�S�'>�FD��6D��?U��5��Z�H%\��-9�>��hK��q�N���w��=�5�E���S�g\�
F�9�e�"#`�B��.	����ی���1p�2�lj��S�yi��=^�#cYڔ���§h��D���Jƻ��P	s���4���$�,Ž ��QK@,�e<o��S5�ӄ/�&��w�+'��!�ًD
z���Ʊ�;�tQ��s}t�V���I����s8�PK�D��D�8z*G�$�|�B~�b0�V��v�s5��%��vض"�m{�:�2o�I��y����҈	�B�5Q�;i�N��c�����|�ǿ�a�FF����t+��yv�?�2�~^+����b��`��{ Y8���'�5K�6�϶�{�*Q�?�eE|�}Ϟ�H��w���*|�|j_Y�!;��97⧤|�5�砟����)�Қ�����������B��t�9;)!��H�Qp��'��p��<DMe���N��3�W2]�|N��h\��� ԋZM��G�1�0��t�='�e� �i�3��`-�����!�=$�
'��y� �+v����j��Ot�2Y&"+�H=X�P_+=c7(>�V��b�r�-�.1���V�-<�	���[���,���l�`�WAƥ=�����ͽv���6@���P�޽n͙Vu+���P�I̞z�^͓��l�'��p�5��2�?X��o���i���%�N�����셴wI1�/���~��m}X	w���v�4�yP��j�l����8�z�7ͦ�mfdn����	����K�h�n�R���n�r_���}��C�_'ٖ!��Z��D�.�S�F�d̝�wL(z-߰�@!3*Z��ؐ8�;p�w�������ʌT���G۩�S�l�21��q��[��
�c�1���Es��R#~���.�6S#
��	�����B�BG��!���I5+|r�����K~v3s���~���0z����ޚ� ������
Dk�[X���q��>�/z���i��&S��u��,���'i�1a�,3^�N�هLV������|�!�i7⭿���s�`�th.x��,���j@�.���p���o.<J]T(TN�*�W.b%m@�"H	��`�}�^�g>eO�1�C杄�-�|���M����!�Kڢ��}�<Md�����`�1j�ក¤�7IxY�qn��^�L=V��AR�����7�e�8<OG�� �Hhi4������KNE��iY���?�wa'8��/(b��.r���13 O�/5��^~H �^v/��7 ���K(ЅWmЊH+(16�ۨ1O��g#��!���ǌ@wG�Rm����臇���}D��?�ad�Ą�r��}+>��IBi�Wv���⥹�B7�ؘ(�m���>и���v]�h=��Ё���|Jd��R�0���s!&��xE.�n�A�t(���DMLd�d���O=�?�Ƕ������t:���0����iU�v�M����S,��5��$��!�OP^ڢ�u���=uPgOl㿊���h-��W���������9gq�� 8&�gj�ű��^K�@W��[:{�d_�[)��wm�_�}Ł��k9��^>��	�˂��4	���8�=��լ�W#�%mb`T�����bY<"�|W���z& ����O��MZ.J餚n�tw<'��ݘGެ�z�_0�*),��E�]s�����Z�����'e������2�m��au�?W����t#D�Ƨ����f B��(�\�	N��P��X��\<�%���c uy������p�XG�jQ�ɶ��N����ew�IB
�t~�D���0�)j9<F�:B��lԂm/�e��gH��w�o�g�n�n"i���]~���-m�L:C����K�.�DH��rq>�B;�vdHm49X5=� �z����ҳ"���w�'NFb�	y\#�%q �\������ PR�x��4X�&���X��)ު�gvL+�6�H�
���A��)I�q7�@�����QXZ����Nʛܲ�:�y��W����B�*��
I�Fo0�����(_M2�*�Gx��ų��F����6ؕʹ��f>dH��$�"]�|�q�>�Z������n���"��#i9�Ĉ]������{�]J
�b�C$�b�\a�ht׌گe �8�/_(���O0�i
}�}�>���T���S���\I�#�������߉�p��Q��P���?) ����{g'/�x��(4�Z�c���/^��L0TF��U�"��=a]5㞶@�׼|����o�������������`���狃��,��w�8� �a�������ͤR����g�7�a��ΆV����E��g�J����yģ-�@v?k(u*��P���a�>u�ĹK�U/�T:i�p�`�n&+��L8W�Q�?��S����wu�RG�4k2'ҿ2�����E>oUkVm��"R��T�-d�i���.���p_�&�
��ͮ�Á��L�`�A�|>��WZ慴ڷ��Po=��ˊȧ�!N��t3��m�|k�I��$0�J͟���'w�b̷���3NW��ӆ2��ޏ�#I�ły�b�RP�$��˙�:��,���\CA��漒w������*���;���U`5R�/�=dJJC������q�"`��z /��'8TObd�=�"��C1�e8ȼ7�u��#���+'��g����PY�b{���X3ʫ�*��|��� ��K*��ѯ~� �Dj�d�*������4��dl2\Mכ�@�ڮv�.�E,�Vn%��X5�.�6OD�d�L��D��J0�7M�ڒ��(ǄO޽�#��dد����U�>��Vؒ�������J�k���ar��s�N�
kyi�D 8�I?:[%�%�!�{iPm�Z4����+	1�gc��|��}>tg�̄qlqA��/� �t�p�&�MFRL'oƔ�uc���4|V�x������$�vl�J�$���YO8B��t&�W�^3��7�c����"�&�)ԇ_v2�w>��VC*^��M)a�#ep�ܙ-��fd���w�x'��T��05�����>�w\�i̦�j/��`����Y�=/!�UQE��M�J,��Q�o�9T�H���E,~�,������I��z�JM(H0�mi��� �N�;����5h�cq}��t}�w����A�2�v�YvWG��v�<���8���p�Aľ����X�b���F���c���3��P�����C����	��'Y�Tr�#���He����!^�7ٴ�Ǽ��yl�T��ߞ_�F��_��^�h���c�&��������a����������՘��IQ	Г���Ny�F1�	
N�`����G���,Y_*�%[Ǔa.�[��u�=���[�+�u����F��ǐ�d���w��Ŷ.�X���Z��s.|NP�{3O@�g��ݰo�E8�ʤn�gV��=����#���:w�R~r���"b�a��"Đ`��Q��`e7\�7��'g/��>!��]��Y1��Gf�a��|Q-�������o\�Vљ3�umR�K�F��3�ͦqSl>O����1p�2�n���w!�9a��2Sv�m��g��2�f��֍DO�sa�Y���c��yv�ݻ��UZ��f��:y:����,��,�%��rx�Q��re����)Ub��&�Q����>bN�&��p��ࠡ^z��V0�h�E<��m��yn��L<?^�,XX�B��>9O��{C=	bĔq�6�z������]3�r�UN5\E8D�2�ӻ6S�QH=�߰�����m ��'%h�{G�Ά���xE?	J��57���^z��ک�I���c.��zކ�sz��9J*���E8a��1�͎ҳ���l�Z�R��
��ј��%|�j~����qG(a�0�S��D3ܗ��Xzv�J��+W��뭐��+UPJ$��^#����]�t����?IŖ�����fvy��L����hX:�5���{�Ǉ� �8kg*���S7�D9�H��#�ݾB�k��%f�2�̤��s���d��޹�Oqlk	fU�i�k�ڹ��ZnC49^[�5?8Ȥ��� �u����@ǒ����2)4t|w'.��L1Ä�I���={�G��C`�ws��b�Cc�ΡQ�C�t�4�C`��q��wQ8��i��%�?���n��Jmw�DQ��4S�	��.���ܛM�~	.���;'_���ۿ��g���v�/���O�
�c��E��{���78����y��#�s��P9�!I�1�=716I)Q���}xH9�W%T��[�w?�o�q����P�,�7Ov��I�okr��L�a�~���;v%�<uh.���Uʺ�.�,-�`4�l�L6Em�l�T�2��i��g9��߬`ţ�R9�Y��D��A���paI���`cE�|,"���w���ϩ�?w�U��ws�λ�tX9g{yޙ3����"J@��0�Ϫ�X$���$.g�^'9?�������������&�I�\>;��U�at����@������~����ƅ�9�]˄�-U�+�oGHPQ�ԜU�9-���n ����CC��h6S����2Ǻ@�Fo;�bܫt������gB��� ���r[!L�y��p�D�>�ͧ˦�5�Ve����WTfsW����/��o�(3��DG�o�:˓��9QU>�+D�Neȵ��/��n����dh��2Lv��f��u�bb>����-�ƫO� ��l/J��owm�D���:\{����z��*ʲ�Ih\`E3w�a&"z7r%�1�8�x��	l⫬]�f[9��:B��d��z��E	��h��[�9�O��������qb�
��;W��n��z�f�ꩰv�7lC��̩��S�@�kOxp�_l�\,j�����t��R�J8�؈�S�9�;h#&��Zb��F]R��y�?�:dJ؟8���,��f�+�"������SWIXR�f�+����-�>eI�&PդG�b���|V_ڶ������ͤ]�p����n��MVW~�&�[�}}���2�%B�A�X���5j�^��A����-Lq�������W�D��ct\l�����~l@�~��<Vd->y� ?���(���4���'N����#���������-�rb��F�h��z��1�3�2�==�D���(�Ve��˘��>(��k0�����(�o����m�uZ�!�<�:H3O��c��{jh)�d?@�Gu�*b��f"��I�7�D��� ��5�T/W�#�C��(�L5�Oi{��A�`7X�hN`4�0�B6�~LOp���hЃ�f��)r�mt��I�;�R���/�,�D���#��ϝ7ȒY���+f�~�V�K!]g��4�`�kǱ�=+%���G�����o`�Y��b�k���(ʾ���� 'nr+H���ѴHLb��u�<�[�G�1E�t�`�>�t�{ՙ ��H(e����i~�.���ś�-������p#TD��YA]H�N�C�ݠ�pPA�^`jO1ol�����(���f6��Rxݡ'���&As]E�Y=��=�[�ƍ�S#{@�����ْ�q�M�ѣ�E�-�^��L BL�)[[�����H���ڊ�ѓ�4��=��v���R��57�d'�W#�9���ء��m���֐��0��
�pZ`�3����
f�Ե�D� ^�v�Q)�Pە�>2*X�+yc�JKU���Ω�D)7�
	��S��?���p��R�R1�V)sc����0�����SHs�KN�G�y�NM�~�ɣ�[�E��=��Z�؛�1-�X��e���0�C����С�!���Q[�(�[�ȥ�f�o��	#&��N��'�s+�cb����L:u����x��Rc�_*�&#��)�����kv1���>������u:5.�ŏ�i���M����<v�q����(��<�^�p��!+v��%Α�6���j��D�ڀ!&�ǟ��jv\x}R����7A~iP�}�Ċ�,g�!����	7;�̖aO���c�������C�h��D-g��&
:�-�"��>rҭF��Z���wZ�O����<*��:�8?�9��`m�-��[NҾu��f~�^�י#�y�OjZ�,�1��`��� Ηm��75j}�Y�P:�G=�2��a�*t�E	�֦\Lrx��nKv���g_y.�=�dv/���P��˵ZU�}��-ڳ�S_Zk�F��4qÙ�J�I�#C�b�_�,������ǟ�v�H��v�N�*�٧�w����?�)k�1 Dl���"��c�[�\b�w����p��4�U�sYx������m�#�?{䄫�������󕴈��� �qn�W|�߃���'�����|�b܉[�#�������vy'�i�Js4�}�%,�2�$�2��F��b��D��ύr�)g�c(y
1�/J�5�v|��;^	W�!��wgˏ�n���Zd� �v�Ġ����J39���z	��a	����)�n%����������i�ːi?=�Oa[�6XS/�|�Rn�EK�;�+m5I�b܌ٺ����U�����g���+n�ܑ7zi��f��TC� p<e���X\�>�9ll�:T�X��lBi�r��j<��B v�eo�j7�t�/�E\�d�O�|�f�ϕ���f�=3����$9>�dE��-*�B6�ԏ�w��y�`]r>7�ẨS��A���-$��ɫ��М��k�2�����ӧ��]Z�CP�9��MDp��<���9+�N��"t�$��t��`D��d~&t*���ɿ�s1J멧��M�e��	�4�JG��N��Ο�=�(?�R(82�ϻ5��砳&$�R+ߙ�]yXF�o�/��L�8Ja9i���Ԙ��k�����H�#[3�أW��(��]10�ɺ�-n�'I��UxO��<w��?g�㍊�c�޲��VY�n��ӯ;H����B���ޟ!�+� ��=��c9GΎ������dl���o�|����A~^CE��ҕn@���J��y��*!�N��J�%n�G���&ߝ�!���9]i�b�='}x7��*0�(��Z�N����P`}%����v>���Ƈg��������m4 �WYd�g8H.���{7��A�:-K���d�v���,4��=�)8y��y�bFu�A�&�[��r�8./v9�sЅKzĒ��k?�w�[�����Ca1Ʃ_��o��p�R�[�E�H���g��~��A0���P��پ��&"�NFgz�<U$�4�/�u��B�4��l�>,s=Y�@B+�n��]��<�ڃ�ҏ�����q������"�����
�+�w�.@��f�ו��ko�ڦ�!��i���)ہk3֌[4��&g���k�N�x�F���� �E���W�"�4���YU�����&�7\&l���F����_�Ϊ�ZeQuL�����Y�?��u�;��<���c?�4E�@ʩ��Z�ݠ�K��Y+�@���OXf���C�B�MXM��F[q̓v%��7��('�:���+9�����-+5ˏ���Mr�
J\"�V	蕺����?�:�n��c���!ݣ��P	k[M��]��pS(�A���Q��wƟdm)D���B��kN�yz�6J�6,O�l(�O����F�@Ɯ�Fv�t�@
kғ�T��^0��}��q�2Ֆ������5����Ф�.�p�O�jd�0�8߬�����e��9�t������^���7��g[�G�T)�=��:_�V�+w9Ⱦ���<L5zd�U��~��L/�)_�f��O��JzS�}�qPٜ� ��vWq��ö�J���:�=Xh�E�Ν��%�=��^e)?_bXo���	}]$�͔#"��,߼�"��=qyz`���'��_|�OI�E��4{a�%��-%o���c��C7{6*IB������v\j�s[Wۘh�o�}i�3{L��Z�\5n�"K|��9U,��J%�>�Sn�h�-f�U�mȘ����p��'��m|̣vy�%}{Qٯ�&{�u�x^̊�ſt��&qp���%��q5�����7�����a%�\ǥ�� �Ք��mi������ڰï��=tns�����o�vB���+sݎ_��}�	dh/x��*�s�c;��O��}}�1�#�/9��^��r��ً�*r���B�K��S�,�+0=��hQ-��c��H�zWҾVl2k�M{4�˞��=�Ѧ�D|gH]\em)MB�աG�l3�M�1�At9�ןf�Hv�~X�<2exw��M��[LO�^l�gKX����u���n�챼o��w��*�+)��\/ ��?V�}�^*'���N��Go��`�-��덵��B��b��� Y'瞻; �:�uf�9�|4�*=e.�܍a�Uoβ�E��
��lX��@�.��h�!�11�q� �"^�� ���>�n�^Տ�"�$�n�]��8�XɈ��9.�9�E��y<�o��ߘ�FuqJ����2�;����S����-N��_$'bs��,�����Ɨ�-��ŵ��4�E��m�����g?���XtR���>�K�=PO�>6Ci���n��'륈D+'��1���_XC6�E?�����y5?�ͅb���'��K��0���s��R ��q�o�0J��u�8B��i���׊�1�O��v��i}(��^��3��-�{5'b�q�� ��� :�W�'x�X��[�ց���o�����d�A�}=h�o7�$h�����g'��X�%�A"\|��4<�t�
�gncB&>�Aր�^'~�UNs``/ ~���|9������X9
�jh�)��ӀJrM��ʺt������Ki����
��YNb��X#&dj�yi�R���W��z#*WX�k�f8BM�?�l�~f�V�6��\�p��+x>��r�&��}#�҄+Y�S�F�Tn�-�lb媦�l�M*3�������ݷ
�G�Lj���7�v2���{%.8���mw�����v^������h@�o����p�M���t	_�_��&u�6�_F$���%.!�{��*zG�~�d�3Dz�]�����0S2}��/)���7��DU�Bg@����i���nXE�M�[z�M���i�N�ύ��!~�������[��Hɽ^����6E��n�_(?�z��B�z��Dt~(��(�A��?/�!���WL�A���CV΄�Ʃ�w�+�%"�hE�{В�+�m,�:���ĳA�ڬ̘?'ݶ�dF�[J����h��[��QҶ�g�^cm�����r�� ¬q���;��E��S�JO�%B�R��e7�ݚ�X���P����V� )@P�M�d�ћ�0>j �k&?�h�7F�����-�dMv���UL���ӴU� �F�p%�=-���^˩f�;P�ַ�߼ &�'�_���F��N0L���0-}u��j_�S��[�����=6�c3jO|�huoI%��˄$����f�`�HxR�+^R���V�6rU]H�:��%M�"�+�7���G��v�d���%u?ؼ�8�@�Đ
>�jt���4t��azi�.�����0�I�А,����V�z�+�޼�P��CN̡�L�C���3g�"����9��E�S��FϠ�<zaO�z�nw�ff�\�!����� 1|�`^�Y��M/lxEلk~���<�e�����Y�c\nm�O���w�l���,����t���ic��o�M��^GN{z�]9�[���b���/��h9�r�<lR����ЄZ��lj#�$�AW?�@�b�İ�Cr��cS�*ç���#��Z#4��F������[�a�$1����`G&��;�����S�
> �ͭ-����`�O�����\�
�����)nx�b��u��7�j�Ŭ�T�t�|� �GƊ)[��c�XNBy�>�|>�䐅 V���N<�SD���.�K�����������1�*�����3K�@�=�ڗ��Ć[��G,6b'�����7O7-c���;m$�'�A�x�o����,�M���.韊�>�\�o����O�J��f�U'dؽ�]2��eݧ=��ǯ�`K������]��訐k!������'�f�Sy Ml �uA����K�?C�1�Ѥ��1C�f6"ŏ⁐�":�pZ��W���R�2?*>��D*��Kݾ�����-D��e`�|Z,1�.�^��r+3I���Rǭ�`�+��A�©��k%*�H�/�0sz�y!�D�YlK���1"�7Ow��]�Z+K�� �^�dɲ��>_����iH� ��ʴ��>E�PR�#�M�'��:� �A����b?!��^_��2OO�7�ɛ��+$4�����8pu]���U�? �1j�V�:���0�[f��k������J�u��&"!�d2X^1(�i�y��.��b�,��0!���r���V�^�%c%���-<��j��2�l�h9�;�S����SCe�n���Ԇ�~������ȩŊ�Τui������
&����H-F�S(����čiq��:ιP����Uc�Tla��hμ�!���')��%k��0��W��1�e�f����m����O��h���,�n�\���|ŨT�u�|�
��S�²k��U=�J�����$� ���$M!�?$�YI�������%��I��(��VO���<Ă��7R,f�>�D�GW|���A����7s=l�dP���!T �_�'�4F_�ד��9b�L`N�I�9�����b�l����>�;��s7$�d�UY"�[2�ɡ�����)��XK����$��?���o4�7'��X.�{_�'D���� ����$����K�|�'�K�,�=c'D��jge� ��'�@r�aw� Pru�β�Z=��%+ک
Pϳ��E3�qӖtڏ=�i�/����<�J�z�A%�&��'�Y��;E�2L��#�g��{"]���g��h�~��CS4��ڗo�	�T�і���-<��4��:8�\#���
�opTf,��8.�"�� 0z�u�J\��$����P>���u]�UJ�*����m!ѹ W�c�e���b���.���L�t1ο-@�J�t$ݦ�H%u�Ʈ���&���8V �%����5%����N��l��'��T3��d�M�r�fe��Ϻ#��,�P�{�O�K�Y%z~���犐���9*e�x���u)�Qa������E����[{��Č�xe����j8�mxWav�k�0Qm�#���ty���W�q+p7m>%#���ta�t''l���Κ�b	1p���kV��7k��c]�N�vu��D���q��!�VC��7=.��Yv��̠�#]Z�^h�Ak?J�3N����.-��ۯ�^a|�:�l�����=FÉ��0e�27`�:9�a_�Xİ��p�3����s,�i#!'��� Gm�zڿi�Oc�\`D�@~Khd�x }����Z.��u��8	�<��n�h�8�$�iԮ�6�c	 �w'�n�,,�uE��T���G���1�ɏ���?������6������GFu���^!�����!<�-"`{n�a���������.�����K\���w;A����vI�3�f��~mc�,�'��V~1g��8�sZz/jK��'�m̙`EWX痜�D���\�e�^x9�x�n�F�C9���:̩,F�#r���Ek���6ƹ[��|b��|"�i��o~��V"����Bv9$���Ҧr4��ǉ�.3��8;c�/��/Ļ�}V+�Xz��ak��wTZ�0K���\ކ4����7z��j�oz�H_�i(�)]�+m��L���ko��H�=؂P���x!���[#֩�Y�����ר��T�0�nLA+XUqr?௜�qe��9�ڧ����sz��b�Hj�%����2x����.�=FB�E#�
�O��փd0��V�������Q�~�
�<P����@�2�[�?{��v&G�6Y/��		Ђ��}��_[�z��K�0�<��@�kDr��41��Wbxz1Rn��1�}k_����l@W�0E���ԅ�i9h�l ���'k��P��0rK4�,� ��g����vn�����*�M�S�4��@�3�t������U|�r��_l�3�i$y�#�e�p"פ<�o�O�%�ΎvSij��l7�g���{�c- �Q�
��1X�����[{��v�!�dašZP
�o�Z.O2-R=~ϲ�S9�ǎ���V#G�|ڠQ")��q^�H��^��.��$3'��e
�Z�Xiܜ��b�eF�7&g�5Џ��._�'���Uv/ק(�{M7��c_��/F���+,õ�_��w��B��+�����M*�*�M<����ǵ�w��J�������{��
��G��3��Xw^��b�)78��g\�Dw硕Q*��)=��b�@�.����b�>��H�p�gs8������g�|�Wi���qJ��!�ڨ[o�聇�p���
1]O�&�Q��l�>v���'ɋ3>T>���������1�콘y/���ͦG��gB���J�7��E]�Ԟ��C��]�d�����~���+�67�~���]1��μX� z���l�N�h����9ޗ��0,�=�"���K�ϱ:�c9��n�vk\�d%�w������Ύ������~0 G��/6�7��'���4ҧ�(��k��b�.R��G�@�>,��;츀��L�4��=g���?���Rj���z6'w�"o�&��1cfg�p��Z=��
3��4p��-v�g\D�YǙ))����x|�&?Ž���S�*�L�����`!�-���e
�����=�9�� E��_4u-�'��u�5a2����+�����Y@O��
��Q��G@�Y��0/~E��Zkr���h,|�c�F9!T��-iFӎ|�F�~�Ǿ��d���+!!Y� �5�MR})<�P�2��Z`�;L�I�L��D�x�����OS.}��H������r�;��g�H���p:w�o���=�o��UV���&�,�6���u�d�x�//�Z�V`���:����KS��4��ȹ\?�PS�/�H���a사P�u,SP���Z"|���4��JEc��?Q,�\8���{͖Kj�rF Y%��>����l�}��X4�y��Ä�Y���͑{���q-�]��,���Q S�u@�ݟ��UAX�r �c��$48Z9��݉O��F�ۆ�Ǆ�T��^k[߷<kt �;ϮW�|�gM�.�=o�����!�g�Js����T����@	�jV#Yl�\$Ċ4�*+(��\�S��w�0<�Ih%k/�x�vm�'
$9&�����e�*����+�-@��[i����/4p9+�H�H���ws
�CT��h�����D���hٌ�{�ȈU�щA�D�ެX>	TͫS��Gߙ������L	��VW���/��A\iW���#��(Cw' ���0ù�BF������f�#�.�cR��&�{@}�1&�8(�$	��|�;�Gy,�Ls��y�+uN�r��%�ځ��jSc5�p��+�E���D^�>GLB��3;u���c-�)���p�a.� �E��;~%�2l,u�>F@��QO�2
�����p�r��)�*.�8���r[�bu���/�ؤ�:��I�e����w�-)�BR��a�P�^DG5�xjqsoSǛ}�x�+���*rI��+��,8O6���Bw��d��)��J��`E�he<A)�)7kxZ�,Gp����`�9���"3H�N��53�*3������1劆��/즎�L,"X�l��9�Ư��]�dx����V��<˷C��;I.s�����e^�\������K�z}i���,�N��l����9�݁O���m�e�]C4qKٔg�껪l�}��i#�4�i����c��&��d@uu�{����i�^��
���˲�k�aM}gr��$&��k�v� ����zq}&�\�۾o(����Q�:�ZoL�(h��U�ƶ
��!�f
�����ʛ3�6ǎ������� �P8+���)�"�����H:�-��GmI_�v��̎�|�߃�`�9jL��d�d�x��~��������?�r�`/��(��zM���2�|�����h���\ �!���0�f��oM��1�/D/�.<@����(��$�H�҈��28	��)>�ȆG5=���O�2�	:���H��Ar�wxû�<�>�ׂv��H�=�S>z�����y?�Se|+���tO�1T��c����_j����!ʢP�������{�x�E��;Ɂ4E�0&�ǣ��z�j|m�^��t$�Hd/s�����t��o�S��R=>D�3�<p����5�^�����j�\!����0%3�@��+�%����ln�&�����z8D\:R�Ϳ���2:G��tSӤ���܆�IwǢ���!G�4�	���4�S0�[��_�����xͿvP{����,�1:�%�h�C����?"�������Ζ�4vF��=fmK/p���M�5m��.`����i`�W�W������F^��Ε��a]Wo'4�N��:w�;��Y_K?G�s&��]*�%xf����>���P�U�%�^�|��5�Hh����*/�I2�9z��e��qW#c�{Tb�µ����kB��j��pS�[?��1\* �\p�]������޸��1��~�ir�Z�,l+L�Ye�x?�b�z*��i�P��j���Wl57��i���	%s�ћ��Ji��Y�&�48�"�$���1�MBJ�TDA[�YF�|�8�{��W��s�`x2'�,��V�9`�(_i�v�¢����>��_ZR��Ś,�n��{�Pms �{�U���F�p��j8\h�R�.�2��w��\=��"���	�B��l!h�?��<�}M�*���+���sኮ:�2-�s�#��ϱ{��aǌsEX�(\	�P�E�\�5k�}�y���?�_b���	3�
l��b���=�N���]��FX� d�F�;-�w�Q���D+��[Z���E�3�E���}ا�RE��kV���T�nx~��c-�\�ӣ�0�]�pE"����^�7��Ӷ��a�b>�{���rR�C'-�2��FN2rD�J����oW�x�i����&jpv۴T��'��7��>UR��m`��T��8���8m���Ɍ�cC�q��w�W7�-��U����Y���L/�։G�ͽ �ld�}f���sE�C��Iڕf����8U���4� \��P�?1{��Nr��KC8ƣg�����+g��K�
*A/�oWky�{g~2	�}�`�E{��Dm�͐�݇���=Y�%էy�����[�˲������r�A�wo`����[9{U��J�'4z�~۲=�k�%�Ok�zQ."�:ʇ#�E�2����ǷؤҾf�ܷ��F|VL��\p+���U��x���f�C�|��V����sD����@����j��`����"�~OŸ�98����!�/6s�U���뉅��{��X�x��e�0���m����*D��/���5�'�*���,���u���?���t����u�]���g4`aR��{X���$b�St�*��wMGN5���>��N��p�z�.cZ~4oȮ���k�t=�{���w�VxxS���d�C+�7�3v;�G
m9��׮�[@���tnĿ�2��23G�1kO
���(>��m��SE�l��iK�+������i���u��0k
�8@<$���%����t���\*��/C��P?r�����F��$n���u`�o���lHU3cD��r�Y��n�����:��H(|�a�`AIy��7o���c�&d�� |�����췇b�hbAT��dIG����K{�0�����tk}�N�4��� ��xHˢ�<O����7�~�*�w��w�*@8
4R*�`F�ˣ'�-�W�s��98���R'���{��\����l��S�ǹs��A����Z��l��JVOo�۽C�C>�
���q���,-�L���5#}�<GXk�<�|	�� �����zb�^�6�n!>?���YL%J�� ,�ة;��\m���A�H�dt�i�MDCqј�}���gzA��S���2:cL���ŕ ��?mPbnD�`���J�'nQ49����,F�XOi,Lz}��-lBǍo�E�����E���4ھW����{T���-�o�e7��W$��2��P/(qTW�L'U�%p�R����кL!`��o�'.�wC<G�e+$J1�6/��z��mȽ�I;��{Ӝ"[H�� ��L��k���8���.�1�GHZ�4�u��k���K�;��
(�ۼ/k��z��#��0Z�*�����vu��r�
�d{��1دJ��떞N_�&��Q�L�7����Gv�3�O��=����2�k!ٚp^:yM�?m��"LzTM�En�`V�������X�V�%<_��&(o0��"rf��Wt�D�;�<����F�����m�л����ևZ_n��w���s�j����a"�'b�V ����A�Q��!�%�Z� 26둥ow��e(�m��@�p��9�Z����D�
Js�m�G[J�p��q�2������(��YS�6�G3�]��A��Y���&0j�gI ᝮ�	��w̔x=B�55��E� I��ݭ�Ϟ��
tȷp��B�8���ۚ����oX'�c��wPD�}������r�~T�D&<9�;ihR������פ�!�J�,��suǏ�V��H�@%!��	����ti�R���O�3P�Y1pC��Ԋo���K	��R���pD{/��S$��2�4U�$p�Q��
������ǉ+�V������:l�]�9���o�������*Ң�u��P���:߶�_���p\J�>�����b��ͪ�$ ��vԎ~׼�4͠�������3���'j����6�h�-�:�#�0��IP�<ǥΣ���pF�DYoI:&B�<���cclك��i���%�s�K ^��-i�#;E��-HM���<$-���muW�W� ��+���	��'�S�5��ņ�H��!��c�QI�����״KjF�G8�+�� ��ŧS�񝺧���MOr��k��wKn�ap�+���w�FXO�_��qX��Oc�zj._�:\{<��h�:v��ļ�3��dh�8��Q��H�}�^��tv��;���׺��ȧ�ȝ��V�	��H��������y�I��H�-�����2.�w�ϖCz?O(Ӌ��Iq��2�&�U<�� z�Y�)� �-r�V�b��-�Q�<B�..�8��NU��##r%	�l&1>Gm�@�Sv�;~���et�l@���tG�x$��{sT�{��J�{ɼuV�� [)�-\ \�7!o@s,i�KOˁt�+����N5�ŧf '5R��������Ǿ�'Ԟ���+GT��]H��N�A&�����p +�T�"���>�V��aֺ�.�O�����8��qO����(�sY������g1���%��f� �0bU>���!�kk��*dk������vğ	x������v½��s6]0#��@���/Wm'�_��Ya�Zn c[0�T�*;�%��2�(�YF���8&͔�nk����� ��*+3.��j��K�#��L`�z���Ղ�w$�"n��_���A����$�guN��s^Te �|����G�7��;S�v�D��"�a��,�et����Ȣ���a��%W�2�)�M�]k<{�T2�#K����连���w�Ѷ�YI�J�(�A9������\PH���S\���Z[�s�kk<��F��O�G�de~δ�)��Cy��^_��vY%>D�ݰ�I�|(��R\���״�w���@�����ߺ����zҪ=RYKM����y��ɣ��9*�]�ۡ�u���#�7�}��{�}���*(����s�g��s72k��LW� �:j���E��E���I�4��!hV�� �ٳ<\�|��0���K�����zD��֚��a�}�͙�7-�wREm��cKq�,�la&�8�`��L )��Q+Ͼ<���nxBM�P�f���|?�d ΋�	���ˎ�w�.z����p��"�wF����)6!�9K4�O�����Z��p�`��9��B}%鑦�m���k���IR�]>��q9�9��Y9�<��(G�i^�'�n\��Z�8B;�u #^�j�9�-�$T��5[��:�
-���-:c���`z�i�f��S�N���V��`.em�,cK�Xk�#�,'OҰ���V-�5����_�ѫ��*��PbG��Y,���./8�IR��|(�����U�M�.R�<��{l�b��T�jIa-ɪ�'f��^|����B�,=z�\T ��۽����Tê=oT�/!��RVV�[�+����)����q���P�e$o�F��rܫ����-��6���b�Q��}�:�m/�l���m=���&a��G^�� 萢W����Hڳ �Wv�f���e�$�ȍ�_�K������{��R�`Ȼ�G"�� oqf�3P�_�z��mG�'���X�@���2㟠�u�����ɦU$s�}zwGq6��z�#�L�t"ջG�p{��H̄�I}�u��_��/~+eI��B/�3�-��l��tiG4�&R���6�G3��惐f�B;��~Y�gHcc�A�q�"�%
��e���
S}q��"5�$���-���uw��#��"ru��uF�,/7����¹0���U�ѣ(�+mC_�E��Y�
�i�fY�:&���y��Q���w�?c��1;Y���x'��A6O����U,R@Z1�A�5�l@#-̿���^�{�b�?'&�eȢP��L��N���+�V�-��I�ð�/�2 ����O�mq����,�Z��q�K��V&穸��:g��q�
��w8%��C (P�V��"[�o���G���X��#R����x�l(���x}{���;��W��*�P�Td�R��ś�>�C�qD���
�Mj�Y����]��4��:�4��;}�:�_>j�g쭬J��̰X���NT�	T�oex�&pDg�� �Yu'c1�,�
��j����(I���O�G
�N��ap�m
M���0���
���);k�ܤ_[S>/���1z��ez�f�;�Z� 	�؛��ӁI����l[lk�=G�߆�(lI����pE�#�z������r$:)6ZO�jT���oڵϐ ��
R�j�@��H���$�4?���%��_�;�[&����Y��8�L��.Ȁ6a9�.�.�H��S�������5{�<,:��+�nM�i�5�k��\.j�}Ǵ7o�O���%�m����6bt���9��%�;#�Q���:�*�,H��/HH���簵�{�b@�,Q�P?�����3|����e�7���豢��� d��	������<m��=�\����Ů�E�N���.Xԙ^Jh�-
qֲӞ�	�J2sf1f��J�A��� ;t�2@�\�w�M��;~�Ϧ�U��P� ��w�*?8ba�В\��o7B�3S�rwG���=F�9�[���vs��v�7����Zm] ���N�bTT?�p0��ݼdj�.3��d�L�B����|:9���<��K��0j�AJ�y��/��]G�.�j��I��F7�LqDn��P�eü�4O)��N����8�聭�C<��KDUHt���� �r�6�����lw����HNؒ���L�Y�xu����0?����Kr����_�SF���;���'�ΎWR\|_6�H������
�3�-ӈq���<�1��_-7]m/���մ]�&�EyL�Nߝ���ܰÛ+182$d?�W��$��B�ЋfD�AXMݙ����ѻ��|�cJ���w��d��(�u�������IsA�y����G���P읋��)�L^�8g�_��^7����V6�K�Ӗ'��j}�)�0U	C�t�U���L[���n�=Rz��@ڴ�R�"AϞk�[a#o��6nm���I�hq�	�G�3��Vg���W���n:b���	�x��-����"�]�{�����顯k(�أ����Qмq���#a+Ô�# 3h&�i���a������P"��y�j63��o���5�F��
�r��`���n���M-�l��x�V��<�%�Fp=�����J����~�wNߎ�`�t��'�F�k!`ɧ�����]�䜣L���?θ%R��r��ʉ���(��ɀu �/�*Օ��߭�C�KV�����G���`�o&QA]���f!�_��9���j�?N��:B��uOw���7Џ��;��EJP��B*�fS�9Vl�?9Oj@���K>I$aw%��I\��Z�$9�[뭒䨞�d
�����p"��|�Hy�,5c:�%�2>8���Ǡ���=��/�.�~��{c�����Җ�cCj�Ш��"ST<�ꍣ�>�)<��� X+�wf?�L�m����@N1�����9}�$��=,i�4�YȆ�Й��፩���������8��y1���{�ׄg���3"|�,潀ٗ�R'��%�s�}������K]���.���9	1�U�o��),������E|�Sy������B�,��!�i�:�!,l~���di��J���/�k���C�l�J���.7{5:/�w�O��E�%��#�dUlN�I�+�$��vlU_	��	e�Z�v
�-�¸,{�d�{��5:nth��F��E�C��M�0PUBl�%����������Z�;�>[�A�$U���Kt/j޾(�UŢN�.�z���H�46	�k*�V��\\��:�
a�J���W�1��l���S�Ĭ���,>��
�B��`8�����Ł�8���y�J 9jFN���Y�Z���3����y*�0�U �X���T�1���џ7�7=96���v���_cAq�`�kP*�n�~)%~u��c��m37��c�б]h�v�2>d<%��:_�l�t�O5���{ ��P�ȸ������K`��,�~z����.B���#��Đ ��"�wOGo&+��FXۣ
�;���=E�C�o2�F����4���LS������-���0��i�+>���@�#�N[���Zt3���C��$�?��n��E���R�Sf�wu=�����ǋY�%U���9��q+1U9�.��u�z~���_ĳ��yYi�߽#��o������WUV�\]�M'�h�GfA���R�!���Hڰ�ё��s�طDS1�!i����g�jH%���X�h�ϯ1��[W^�
��i���l�* �4�ǒ��Ț��������ٍ&a�
�Z?~��9UI\}�#����3w�3f;T2���(��F> "�t�/3�7*G�}���4r���N�E
�Ot��#E�(�L,�8�l�>�ΠL_I��.��@��F"	(���͇pގ,����j�o��fS� 
�Yf=��>{�y�����[�ݟ�T�e��A�f�l�x���CکF��c�͈�5��7?��@��>��T&��Na,��'C��b��j�yt��{5�pPK��Ն�����֒��R�"��,��.��d2�C!E��󫊚�On�Dd�g�z��/Cvy��
��z�����*ǒ�� ׫-!Sճ��/Lo{fb��E�\�x�4ur�mfL������3�!�m����'nK�i���1��w��?�E�%����:Vև�d��t�+�E��#�5:��Vx��6W�<؞�Er�u�X��y�|�W�l!���#ė����y�ڈ!@��y\�=&�W�F�f�����N��|�(���s�&B������P�8���&͛�B=�0�	��;P'f|�<��_��E��'���}�n8��Ti��5�P�%q�Z���EeL��2eF1�2r��y����Q[���ڬ�4?��]�)��Ҧ���!�_}��h��]b	k��ޮ��-���"#��K�xg���Po'a�o5���{�J�[*��@�[�wV�K��ݐNP��QR���>I�,!�p@��Ѻ{ �U�]
L"���B�i�zT8��.�)������Uk�r(�����b�_o����\:�K� ���}���,.�
�ɍq;�����:X�m��Ps�+~'�����_�֗±W����g��9�L8�B�~e����'L�l�CZ�
�z�����s�V�P<�}��K�ΜA�%划*�7�v��Vq��)���l�4AAorQ�R�>���Z}�?��AC&��d����N�K̖vJ�lkPz�$c�=Kkf��!���t׀�� ?DD?�N���:�zÑ���Qd؂����4�4�|�dpQPP��Q�V���dhtpRک���o��a������mb��fQ����.@��'Q�<y��\������C�>�.vAOY���E����g!������Ȼc�/������!�F�4�����4 ��6�d�4��
��L{��^̇���5ܙh�r�w쵻O�)���e�my@��((f�z�HA�K}���1�u�H��3Y&[���m����0e���.a?�m��"��b>1���E�C4�eTc�
ѧ�\�Z�&��s��	d��H�e�$y3�ڳ��b�-����,�=��.�a��z5�'�C)MH�t�E瓃6�jkM�P�?�w$�.�㔬�c�o&���s�9	+:L�|GqC�G����ϩK�(��^;��-��9ug�kR�&\�,���$o���|�Vs�F��F����fPV�L
���u_�&9(]�>.1Ӈl��&�.��G���ws�H����\EG'R�I4�ֶ����۰'��0˴b�N�′��zyj�+e�g��c��yǰ�����L+D�;����S�[аo����S��Г_}����5�W($���n�8Vٖ�[��sj�Q�	���*����U�?�;��a�^�.݉�M�
�i�s��㣄LL{��n7R��֞��:PGL��%��	���K�R�B1R��Eޢ�O5�X܀�Q	��n�%>�|ݩ��s����:���#������#�,��Y)�c�� q�ePt*V�M��7��Ђsz���؎���@�C6�s���y�r�P/d`����%M��z�R�t*�vlp�CVX)ܹń���^
������OLm"_��Y���<d�;|ߤ�8_
w�"H-;�L.JV8�bnl�=U$����n�f|�ZU�ߔ)l�W�*�^�#Gjߨ�u�¼���D����J����8Wl%�u{m�^���s�H��2��/�!����S�8��	MK��u�� �rS^u�dy�J�L��˚�yg���혈��'��2��8G�*��x��[N���1I]9ui8�5]���̩�<��d�X�.k��xMg�x��Z;k��g��+H@��:�vV-��<Ut��	�.A�F4��Z6D��Q&����8��糷˯r� m�l�ZB�O>y4�;c<!C���(�z�������t��-4�ܒ�1���l����Bp>^���u�czn��av�Z�{*h���}��X�����L��,?�K �xɪ���%���n[��	,��A��>S�� s�+6>����~~N��l���t<
��aқ�a���yjPKf[|����eM1�q��
2�� �*���F�O
�]�h����\�BS}�8��G���J+�ן��������`����2[$�X�3�f>�����L���� �?���*�D��G���)gt/*�-�-���$�,ߙո�>�g�����AQ~)}�׍"��������b�) ��9`Wc�l���&Pe� �HG���ʬS#�?ʲӵfF�O0w�6T�we�3է���F�}D�
� L��Q�!r����20tm���H����6M쒟�(JA��߻qŹd�f$�W�K��;��qʚjKҠ��+�pL�s�rZh�]�<PG�B���xR�v�m�B�R��o�vFư���k#�"�2/GV{<���H�=k�h�����Wc�NF'`�ن��:6�睻2ԕ����i�N�}��kq\��VN���֕|Er�� #K\H��C�]�!Eb���2��� kbO�R�[�8��ZM������d����jg�/{C+-��p����M����x�8��y$�נ{<����y��PgK9=��b��e�hc�,R�]M�ᗮ<��	MI8���\,{$���Q�@�e����ʋ*`慼^�C���<_�ay��)��K�@#a'��ਕ������x	��j�'@���������[Ry�{���i\0�.���`C(^�VB������o�͖�H\�4Q��n,_jZP-j��e���?fi�H���4%�dǔEL����������3�U���ŀ��l�n$��kaOQ�,�_���9�՛n�b�1;�	��)�k��G�R�x���ޗlcՏ+>��ǵ�f2JߴU�}HlYgS��n�VK�PDsNy	r�t���%ˉ�"�6�����4K����N����$�ܸ3HQ�/D���;%�A�;�i���p,���G�p�H�[��x3��]N�[��<��jG��ϬAb�JB�a�:7�Ǐn$
�n���b��\	D�����\��g�hC�"f"�D{wc�k���=Bf�WO[�9�r���[�-��#�=�17{���H�]sg���;�x>��֛K��(����Z�ˣ7��6CD��Mk�b"f�ࡵ�=�a=J�N�UHP�,
iN=�������/��aut��pӵ��PdMi$����.��F��} �M��T֔��;�Û'PS��2���9?����z��u��1u��V��f����}�T"n>�)�I�yW��+�kn;�^����\�~�j������&��x�^[�r-��[N*ΝPl�')�frv��P#���Y�!K豋|,2�~�/��Ȏvѐ9�'䃦AS�a�L&X��cǜ�q*h®T�H���]�u�4�ay��z�s������.�*-�G&Ц��Lr�C�x�]�$j���U���o��b�Z$Z�%M��R�6UX-�rnM[��,��$F��ɍl�p"&�8�_��>���+����Vv���Jg��yH�B�jՁ������������<D��V�'�=/���� �XŚ�;K?�"�[�7��a0m�q���R7�(���(�4�ؘV��w�U���Wt�1a`Ƃ�KƮ�B�D��Gbнl���'���5'BG��U5�D�Ïh#"B~�����|���!ΰ?m�6��%�`�tQ�ZW񤘠9�3Sc�Y5�#��C2%�\��I"˩�ۓ̉`��Y&k��l[4r�-������t0� ~��F�fw<�4��ϙ"k��Tx�}���*�J6�[?	C�ԜX�ý��ؒ�Q�5����"����; �ɦ�eK���FSԜ�2�l^�h���'i��6�l~���x�{2��9	j�Z$���V"������b���g̜V�.k�ɸ<�؅�����'�P%Gi��?ʡRO[8��K�/L�rJ�_����G���8؏U{*p��Q#�Q�CF�����Ko)��ORg~��)C��:�H'��Zc�e+u���y�.M��8�c1om��eGϰ_�k�lg��n����X��6=�%82�#9�>{�r�u�Ek(�KV�䢕ֶP,�Ƴ�K؍c`�&=�mӍپ���Cq�OÀ�Y��c*��{�:!�u� �����0���'(*����u�/��Ѽ�cj���'�J��L�Tp�մ����6�1�8����>Lg~fg8y4�MʬX�����j_�R_:.G �b�q|��׮W�W�aF�b$����N�jR�Gx��5\��Z9_��4i��'^�,��CJ�H� U!϶�f�d�9�b�qo[5�B��?��aA&y��4`L�9�
�	�{.0�jD2����p� $m���ٹ��F�5l����$Z�h]�`w�\���o+��_R����/��}����A�~k����� ��8Y�Lf�Dcy�'2dFh<9x�e"�Y뛴�R���R�p�Pޤny���?_% c�>����|��k���^Y®\�����}�GV�a�
C<� �5G,�h,��5�ىU�0��R]�6\bФB0�y�2��*@��8�������@�/�{�)����pJ�L��E&/���8�mҖ�tȁ ���	NN �3������'-��3���6�&�'o��S�C(�cݽ0��!d�M� V�b�3z��@��6?����BF�I��T�"%\B��t�I~��1"�^�"���~믲)
���s]Gu �G�s4�Q,����,��@���G����@e��W�Π:��d^`~�3s{���yL$�aQ����V��,r��:�,�"O�pr-Ȝ'����r�+���yG+�����B��Ċ��.��ю5�G�����}a-��vA��]�}!�n6bo�D� �HСp��^�����C4���}�?�5U�����g|7����Ğ��h���!ՑW�AK64A�&a�Rl���Y�΅�������"袬����W�s��8�/�9~R/+4^#��aK.$�%��{|/鵷r� �G����a� �.1�P9�e�(����EP�� ?o����ӔUO 5F�	��/�>)��=D���Jܥ9{~\ ��s��	��!�sf��#��$P1L�A�ȁ�˭[���CI��װ�+yΥ�jBE&%�Է��V戰}��t�{��o+
��1��G���<4���L��Z�6y=��Ю %y��[�q%�'�i�/��|�bG �Z�vs�]=���M"��Hm�ٲ�TYBA�v70�RҴ(7q9�O�_�;�85�S��Ek��Y�k�<����,h���=�.H߻J���qO9��������mSk>�o=��ۨf2�.=XK���IǔV�p�5�~�'zhrS |��m-��6Xy*J��Im�I����9L���hSxx[!.&.���T���Y�H����b �e*�%h�R�?u׻f�れ�_����ik/d��z��5l��іQ�Gڣ���lM���!������?�f��<۸t�O۲��Z8��4;��!�S����VɌϴM��{��\}8qnMX./+��3��q.��� �+1x���!{,@x��+�=>���5	�/�t=�1�=	�+�kOVy����Ó��<��A��K�Pc���&��D	2 �1����M�?���"Ȓ��/Ig�H8�]��o�VV��:e�m?�qa�թ-��B[���o8���=}���R��s���i�(b�kP��������7�A���ϼ���Z;x
���4��r̛��v�	̬��"�G3��l S+��.�N���4n"�)�N��c���Fy ^�:QR����\+�����P��������C�����E����Ry1	��o�"��1`��3�WD�< ����^㎬�R��o�9��D	�>/5g���zԇ����B�"T�kH�O>�.�u�M���R����WT�Ӛ{��&Ff�/�cAk_*�Q��sM"��%E�Y�͙�iB����`UW
G�n�EZ5�5'�'z�����BD���,��:W�տB��П����{b�&�	_���+[C��GI�%�8#v��!��dn?�'�d�y�.���z���3���� �=j�D�F��Ks����YOo[ͻ.B[�Y��o��\[��KH�Py�J�e��Z�����m�bJ� �U�hf �)�2`D���h����;���z�{��\;��n�y]en`�u�\^�L�����x��7�U��S���Ȫ*�L�y>~�c����t��x�=߮��#�lL&	�N�(2�=�8��&�Kx�T���e�yN3RzMM�H���*�3lI�G��	v��'����k����޸�4�<^�=[?.����f�ҍ�A�-3�8��	�`�7��A1��ioR��
lK�0��W�{�v�ylѩl��A�VOLQq�����fpha�*�~�6 �u|#�*�Xb��;)_B�j�e�PE�
c#��ׁ���lʽw.���4���4��>{?w�<�(�yrG�$���`Z=��ג��S��I�nS+q�"�������7*��|"��V�5<�ZL-b�`B91*�}W�{2p}���k̲�&h�օ���u�Ǆ��[&�g�X�7�V$��s��&�x[�[� tCf
�E s�bbM!n=�`R��r�d>�� ��yK��"������k��V�إ��Ax����4��*��dx3�-|D�cSSn�L�U�5@u����g�>�SKA.�hHP�Z����ˍQ�2�r,��i��(�TN�TR����d�8������2-�{_����Y��UX���QTFg|�&��jNHǦ7����ʼm��p��M��e�*�˭g�~�@����5��b����g�wʱ�pvh��|W��|V��O����U�@��Y����z�@ג~���uaI���TK���$���юvVd�B�%�9���S�76����A��E.�r��2�HY	��Y2#� ��-�G^f�;�/��ʩ@�e�'���3���'����ՂX�.�L�)O-�W�^�oCA��Ϗ��	�h��v�2���7Hx��F�V����٭�L>�6����@�"X�񄛞޻��'��탏��2�o>JO��N��&��Mc_�-ƌ��b~to�Nx�E����"<}9����7�xn��8nc{��`�N����s��b.z��U�?�Oq�;���Љ�m�˾]~����{S�*.&il(������S���1.	8�k�{@��u���{oC%���,\iek�Gb[�r�6Ufq���?Pm��{�&,F�y=N�;�Y�xC��W�"�0~X��a�Qi��-���TXx�A��gHc2�M�������9~��OL�%2�tU��������Ͱ����8�ۡg� ���Yn5"�2��1%�r�0��؊��E������e�wH���Uj6�ܐI!�R+�̔���~��a�Z׌@�m�hpə�MY�UZ�Oi5���P�dD�:ga3EL�fp�5�֍B=�6��b��0cZDe>̀���:_�D�ʗie�Oq"g�wO�/�9�R2(��	Oy�wuu��Ԙ^X�'&���Y^ɏ���v�n������˓7>@e �Έzw�,�}��%#	Ӽ�����bN�Վ��	��H`e�L���zڤ��i)��t�'�w��,��a�t`�2�ԺE߱d��p�2Sx%*>��tf�,�"����/��[��?U	�z3�}c9~8QCo����i�zHZ��.ˑdx�����*��r�fR�쁂��b?�뫪�R1qπtLr�.��Yaר���˔t )"jz3�\Pm�EZ܇�-��{�K��]���GF�'��P��hρ���G�;p�v���v�"�����@����q$;��'��U����F��;j]#��Q���{�ron��R��@ ��ߍx4U�r�r�J�=��3x4����}��,{�J�����>���k�������a�[)SVX?��MK���T���H�"�H����I�;����Z�*�G��8�X���x~ې ��]u��+O�]<�9�J}�r��ei�	a�R7����:�y�4�/*�a�n���3�`�9�jA���ol�&bӇ�����ߧ�FIq�UpP�#�y�Z�%k���Q�Nuz����<�)������L�v!8�,����B�$V�����)缹S�|�1��.�q�
��T�]���O����J1%L�.AT�$����E��×+��7�0��#?Ô�B����I�w�=�+*1EZj%oLr��
�v���՜ĉ[&5����Eʡ�������_�U"�v�"<gLUj�����ǶZ��}H��b�9'v��5�D�:��R��z=��+��`�Bw��Ce���[OXD#���0�D��W��<L8��V�\z萇]��:S���E\�~`���c��By�k��7s���{�>����3�@y	C�*!��=.:S=[�/���a
Oy���?V�?>K�_P��߀� �k�����"�e�+�	�ݿ�Ҩ��0�:���M�禋M.�jW�lFr;�$�Lza"��#����Vw	D�"��/��	�Q+Eھ�
Zj䪉���>8g [�>&8�촄��ըGW@:p�Q�� �O9�PF(2.��	^ n�r7��P���~n�x���5�qI�u{�|фDD����
^�����r'�4���ɓ/��X6Gn��#�$���������FX��B�x"��ri*��փ����S��|MCQ��wMg���k�6��\?��T�`[��
H���'1��s�[�Y$|k�\w����H���gj'��*�wLӼ�T>����?�D�U	��CX��hY�.@u/2K�cz@�,�/��e�TaE[������R�0I�nI�����hK%��c�/R8i�����8�橏C)��L"Q���{ծMO|�V[�D���ys������V�U��Ts�W�x�n���;�O�B5 L�#(�J��ó�'*I�Iu���y�wL}w����8���W�ˋf#�BL �Z��W���P�7�_j!��&�aB�@@A���ܙ�PE��k-5�s���t����&�'m�<TZ�P�@Ch�PH�5%D3�ط�d1�@���l�O�P�-a��@έ\��M	�zy�����g�ê���$�x�Κ�g��9f-�o�F����&� �jhN u��G�Tu�s��󛞅P��BN���;?�OBMe�>��g���a|=G_U�bi�!��^�4h�\�6`��q�]��flZ[�1���|��K�U^��㮶� �;F�n�4aZ�:�/��Q��ET�b�5����Ԧ,�`�/L����}>z3��ٷό����A��B&_���eQ��
���F���j8æ��פ��3Ri����� ��Ds��]�͉�5%|V5��V���ݣq�Hì(�bys�� X'B�@<�ٻ|��q�'���"��]%��¾���3�P!���M�����f{ �
�Q��O���gf�f͏S���hYG�U�v,��hjИ�'��;�)q��t�e�6����B�p�'�be�,������|�y� ��.m�,Zu��z���b���I����Җ�������X�S��l�X��a�7�w���,J�����a�T�r�^.�,��*��B� 0�K�eܾF8�E�X�L�:�o�NY-��.��c_i���5훂 c"��᬴S��k?|��9}7Z�?qO�!Վ���ܱ����<'^m땃�ǈJB�\fl�Y޹^����M~N�D䐏dP��:����K�~���w��Q'�������Z�n/[�z��Z9>&Mt,�j�������� I�3��~9ҷ��V�uI�k��IR�￤�VZ����f)��/_`�⛘�W����BJ��]���ny�:��e�܄42��,�|���cMB��,$���2�=�$�'��&���4��۶�뿕����b�uߵv�������,0�%�}"�:6x���)��d4�,D�5K�x��_=���fT�5mN2�V%���K���zN�; l���N&}�� I��Z8C#�-�9Ԏ�����J��2~��J�^���9��n�g &;b�[%EC3}��X�6|���t"_���ąEs]�W4_��h*����>��Ds>�h�`\
qlo�k��!�׬M"q�(;�`�\��/�@�`2JX���ʮ��AEWxJ���qR��K���ym��S������J^1��@��;V��5Y���=�����0<�"Z<uS'�8W骮��oFol���Z��T�;�N��¥︯)6\�f�!e���Ƕ�]�c���*;�U຅g �
�N!֪��{q6�xԿȚ#^(�1�r&�+���ZDq�\����~�spr�4��O,>$4sI��@Q�a ��H(ݴ�c�����Ȳ�f�V��.H1�J���#�bĖA!��*i�~$d@{2z�`�6DU୧�ֻ��K �#`��u�Py���m<�!�#4C�繿VҨ���c�@�l�aU2�]����,F�hz����k�{�Y�i\�e���'�q=oK�8�-�e�-z���u�v27��N�i�4������*W�$j��8W��*<�ePT�2�!BA�x�_ު��R��Z^�z��6U.F畩�
-zjٙ�T（�ǓQ+��9�:�_��s\o��q�ʱO�NWŲ�Y(3h��� q����z7��4n*���Ð���Q^&���y�~��+W��Ϊ|'��bD'�<�\{(t6Z�>�9�ʲEl^��c���Iy�ڇ��:���qGe1�|���=(�Hgρ�ЦE�6߱���z4�}7 b��!f����crg�G�� ���I�K���Y>� ;̰9���ܔՆ�4ޙss!�_T���>N3�q7��
odì��'�םΡ���� �2������ �rQ���ؠ���[�fJR����A�%�'�\�w�wT!9g�],���#�Y�Oط��� xY#�}mģ�]S����B}�a!�c�$��N#�ݵ���֗5�}]^Sκ�Ckz���ž���!�,u� w0���y���r'�-�o9r*�̋�:��u��g��.N�HxZ�M���[��6��q4�K�e���C��oP��w٪ �k��[�]1R��� I��Q�^	�鼔h�J]W-���;vBt`ra���؀cc!��O��C��Vb�'.6��1NӈBM�O��G]�����M�u'�g3)"��3�[B��P�0(�Bx-��2�L|�cޮ6u��U���W���U�����#��m���Q��?�k��SxY���6X��xt����O�>�������h�$���Z��0cA�c�64�xǜ{�=�"�h��;�L�o�>k_D�n�s'�ܭ1��R$VS�������24�}P�����;D��G���I��V�Y���·�M�	�DÐY���G�?��.�f�nXHj�o/j�]c��N UHlH�u�0�Y}�w�d�>�9�ĥ2�5�t��!+^�P�վ�)y��NDn��\���q`�A�Ǫ���P���۽��� 2Iu x�sQ6hڊ���p������D���qy��U�"��S?�z	o�Z��r�/�`VP]�S��Xq���k��&�S��E�M͎+)���"$9f��3��)8�i�ܷp��Q�;b�Ot�ߩK�ߺ�HKϜ�w�X��vS"��b�h� )��a�s.9f|g;�����9Aέ��b�����/�$N�@�k���-��M�@Ƥ"��tR��&�hi����7�J0��4��ݫ����:�8�E�lX����?ݠ���"G�5\��2����D�X|��e�
D����p�Z�,p��o�J9��0�5��]��ѿ�(I��9�U�N���Ĭ,���P�P)������S}h��v0�1�c���keD+��`x�ܛ�I𩪯\xƮx���l���D����S�0I�`S�@��i���2��8����m�r��n��c�=7�da���K�Yf�Q��s��:�3�A7^%�~���)n���"�����P��>x$R��=�oE�g5�]�`�ё�]*�41Aa �@���X'-K��"�!}�d��cmZm��L���	���m����e�X��aK��F�1���Z��/ӹ���MAUn��o�A8
<�3�v�Y��\i�_3M���:'0�QLÎ 1�A��� �R���JƐ���:��?�z�Т�bG~�����Q��A�H����-bL+��6��@��M6[��}�2���(�X�J��`�,�ǣ���q��@�tH:�q��PŚ�?�]��^8����Vm�ar�`�C_/P%�����`��F�}8ɝ�Jd1�����G'>��j>���=^�����q)p#t�)}}��]Ž�4�S�:W��.J'���Y�[�@���$yP!�R��,��Zf��>�7��4���"�#nz8��#\�J���.���T�G �~3r� �����m�"�*�d@�Z�O0��K�O�Y&�������yG�Hl��\�Woʹ<p#�f��Wi!"�֦	���:*l��fui"7igDn�-����+�O�u����gr���и�y�u%x>hS�_-(��m箉w�]���t��.�
��Eq�"Y���`��\���2��(	������G���MJ��Q���>�w�q���#����$������(搻�"��۟8}��gn�ϐ�y��*j$��/gE�g��2��4��1�d�>RY��(�5�1���D�Eߪ��R|�2�T�\-D���&f�������Ǭ�+��Gt���J�^��U�܂�p+��q!�5��'io/������$@�t��v�!<y�S��RŔ^g���YTh'oVB�Ѧ���^����S)�s�sJAuߊ��9tݬ�����Φ������e��J�iB�D�Ï}��3�W�'����5�� ��g���X�v��T)��*9��k�H��ٸ&��o}@j��.��氪�40.t��l��`&�����4Ke���P�<Q�̴�ni`�n�+v��BV�Z�����ݾFos�^���;Սy}��.p���o24p~��+S�X���T?���)�K���-�P`ߋ�4�fq+o#�Kc[{�/�pas*�1���U�#��Xy�'%_���;^�P����~������i��2�^3�΃��ە��o�M'c���}�F}��!�[��ބ���\WL����f ���h����mL]m�\R�$K��:��ae���"X�uX����������]��
r�߬�1b'Bt�=�2'`��(�6,�ϺA�x c�,�=s�#���f|L:�Q��}9x���r3��	ӱ���/�z�fֽI��}��� �W2�E����8U@�Y��1qTw8��=@���%�h�2�	����A��辮�-��t	X=R��W�7�=��&	~��jIr@Z����N��.�f�cr������*+��1�2�?*������3V �x'�N �I�AV:��۠�`�:od��N�E�Zx���ņx��V1��T��}�܅��=r�K:���ӎ��M�t]a��*����g��K��7���V��q�5[���_��c���Y���,RY�,�Au��\]LGT�~Q4�%A� P"_���b�����qWt&m�"���K�s3Ҧ���v��N4��! C�~��_�&����z>,��}���X��F�<N������V!�ը� ��_���TL��m Yͺ5.e+h��ڜ�1��Fl�=�H�R��8|=�;�Cs�6]�Hι�'�9�룣���H�!QoHH�U�a�@�(''ӟ��
�RH�ϑ��Na Yq�ڕ�CW-��4V&���:N�EH��B�9�)Ba�Ma	6��9�rR�E<5�+u�#��ښ{�z�b�� Yfm�#]�u,Z��+՘N�/��r�sh���������k8�Őj<��Q��h�i%�$;��٦��ik?��e޵3c\��_|sL-�*z�jA"*���Ln�:	o��ĸ����j�v���x"l������~�_hPBe|I�)���"�q��n����1�X֬~ Y��CV��5�F�w�s^�ݖ�&���\�a����@�ݿ�"dP}/��jٳwy
N���k)೎\��E�M$�eً\J�#셣��&j4��D8��~2�)�ɖL�^�c�{��BV\j^h�=4��G�<�x�򻿚Q��#>�7j(����*�=Ns6������{�s��x?�J��/�?�1I|繂�U���s��1���Ƀ&�j�Ja�]��p�[��5�ϼ�Y�[>(�t��+��A��)��s�!c���r�f�ձa������}8��u�)V���qZ���Y����N���8c��gG���{���Wa���AR�oL��b/)d�Ty�3@=a���!c�+��<EA
Um����NX�v���6 n��Dub<�jYq�U� ��y�{38���@T9�#�j��0.���۟O�B�	hL'�8���xj3:�۞��JA�Qn+.�o��Xۣ#�{��p)N��Y���\Z� ��P����(��C�d�6fnf��. �S�J�ˆ-Z����6�	�" �TY�I�����2�T�Ùw%TܣQq_���E���yt�����t�����
�����Mθf��~��>��i�:���B$���#}Ǖ��N��ӯdW���o3���Ћ�J�}׏��}�n1l�q���\�3�/�u������On�mY�c�9���v��۩�L*o��p�R˺�Ѐ^K�l�:_�r��Gj��\ %s�>ٻ%!>T���I�t�C`��+S+�i݉���|���}w���nt�3�A~�v��Q%t���� ��ǩU.ʸ׫����%�)Z�]���jn5��h�;Ν 8|7���g�|�}~��-���b��E�P�ZxV���h�$���9D��o�r����U�⸔�VZ�s���,�S�!7+$;v��3?��*F�e=�v�����R�*�e������הV�<�r�0�8�j}
Y�������"�=��+e��^.ˏ	���dl�bq�_�7���L���mWVX>D���l��s�z3��(��"k33O6t�؎n,T�:G��n!�sX��ң�5`�t��&���Mw�Z
�����
��͚�?%�ŀ��"5��"��"�`G���JIl���pz}K�:�I����5+#�Z��'��i�%�c� X?D�����9�=
>�=l7;�!K�����D���UZ�&����E��2 a�P���ϸ�:�U��F^��RQ ����$`�]gj����ֈ����'�R���K��&n$��%{�,��f2�����;;�. E?Y�l��Z���!wZN�)������ib���w��'��[j�`h���rtc۾:�7�,�$R�v����% P[�)��"�wI���м2ҽ�#c��&���
����A�h�0����I&e����Us�ƞr�n"�ߴWC<�/�2�2p�,p��Ly-�N� �� �܀��.��Fs~�s²��~A:Iɀ]��>��:܈V��G&�Oꀺ�,Rn]�MTd�K9�w�|�Ӗ�
�W�#}��t�;5p��y��P݆�	S,!���.�w0�$�)�&��@��Z~�3A8��Jk�t�G<���@�⎲^��J5D����!y���z�q�v�9��'�V�RH�LP;I�&E�1^����Emq'�#q�7�!�N
�J�AY��	�m�5��;�k���������<:�,�gE��<R�(l	~��i���r�s�D�K�����0�	IzT]sd�I_S��UiW��蘛l�؈+m��6dC޺��\Dp����.�'�4�h��r���Nn�|�_�ȶ݀��{h�:�i�e��T�.��JB#�4�&�,�L��@�	�7q��Ժ9�KOl��t�0�#����T�Gz'�ހO6Aj*}{ ��z����\��X#�ˌ_�bv�4`�	sߔ���Kzgj��!��A�qkW';��R~�2�x�W��'���g�$-�N���Lu���\*J���f6�U�r���qZu���{��Uý�]�°Ty�?	^�&�8�����̀�����w������3��o�yA�T^$T- ���� o[�x���8��hʳ�R����$���l��PO���8S8�J$дE��=��qie=oV1f�z��R����mָ�l
�c�u�K�v6�K2a��`�V�����Ma;7j������I��{|e20�k+�������7�}2)L;��WW]�'ǯn�Q���r]hH�qq=�:Iގ�vD��a�Hf?�G��K��Q�g4;p�r~B�L�K �|�%��8iCc�2�U!K��X�#����`*��9�������}�h�/�~��5�i���c�K��[H^���2H+Y~�#A���JT	���-��z�fQ�&�tV��`S�s��-�>�Z]O���f9��j��c�8l!���b�bxO�
���8T4w�D���]�t���H)�é��^�Í��Ť�Q�I)�c����n߲�؉�n,]�:,��Ҭ4�oeT��<�gDMyr��m`en�<3����d5��S���Wսk�d3,���l��v����~��$1���6�0�
��HN�䊦�5�D�ZXH��<-AA�gV �m<�(�n'
IePC��r�Z�5��o���@9�.b	Hj�'����p"��(;�=%s�F"g�
��Ψ*�NQ�x�'V��=�=bL�Q��2fl�9�ӹ��d�w"J���!Q����0��n��	�n�U�Q�KlI�;
@�i�������b��e�kPַ瓣��@=�n�2��(�|c��ʒ����Y����&��q�I���%L-O�7j,X(=(9ŝm���k^}e֏��M���K^f�hG~�1�.2���g���z���|@ \b����9qR��O<���4���������j0t(t�CJ����^o@|��~��4Hkx�K	� ��'�%妺�0\)��K�*�7/��1��w�*AQ% �"��xD������y��89�b��H����~��B�׬P�$��Ժ>�+�9��y'���dkPP�g�4ʃ/uRN��4����o��ϖm�P¯ ��r�,
�[ �C�ʄ �O��iv��N{�����s٭�S������}��kIVO�����x'��C����$X�ܤ�0ы��Y�����z�2�?������J��?�]9�H5��U��.L�lt)[�3CZ�,��F�c����^s�{5_���/.�D��6�&���9o�:�1h�K�Y����mH�>kd^K�2n��;�P�BW�F�\�kj�'×�h����LT)��BO���Z�QX�{'a����
��ȖFz��� ��b�a��dP��I���C(>���be�Qy%5t�cX�K>���� o���!�����wF� �5�a"�-���9�{P�����!���T�-߮�@Z7MC~��G��(f�,!�yӵ`�W��lYf���VE`�����S�Fb��̥��-�ڨ���A� ����YӇ:%�7�1c~����ag�5�Z5k�Mb#-�9���xے�퀉�ß$&���l�=�,�ݕ����:vXz��<p��N=�0~L�x��7Ĥ���� �9��OH�7|�_pƄ����vv�ŏ�O�~W�sf���C�l(�k�fK�e���Xn�Z;��x�F�l K�X���{gOQ�l�8Ž=?�e��!+�sE�]\���F�+h��TZv��e�q�w�c,ֹ5°H��dD7Rao�E:��M�1���$�ԒQ��[R1=ƠE"_��55��%�h�MN� J�Ɨt�	�A˯U�8��E�4)�r"��❷��5�;9T�M�Dw��^kx��Y:C Q�<��!T?o�o2���v ����O(�S)
�K��&�'�i�E�����n:^p��C7��M;g�D(�X�L�Zf�Ss���;���:ԦME�ES�J���������3YJ�IӇ ����ZT��	s]������)��KB��_`�́��%��
HM)	��F�Z2�U�i�p��oR1��x���?@��̫�oJ׿��x���}*4��^���� U�7Y*��#�d��c萕��K�������DG�6�RHX�n���1,>�2��T����;eqPMe�{Y���@oh���E���>W~!�$F=�>9��<�a}a���
���"D�k�7���{K֏�? [MX� 2��8�G�<�ᯫ�%����hI�Z�p�=��c�zA���v�'??�G{�\��Fӑ(������󙽖9B߿�����s��T'�ɕ�j�nspk0���/�H� �\�JZ�.6���z�!YdM@(�L�D�[=6+�*L!�Vp�_���x���y�Z�%���>��c �$t�|=y�-J� 5^fj��qb�5��i,��5����G�-�`�V��iJ���>��MW��|�nAe7`~9!�U�Vd.Ueq���YO_*���i�N�f�S�ė�,�B�ŉ35�߿A�CɮjD��w��F��{�U�sT�WG�:�>L0�wdM,�:yv�^�2��綞����?�hxi6�7^k��ȧ���ʖ�VT6+����LD7�a!���'-��}J����RƂڀ`1���*�{¾P��&՜�h�A�qVc<mN"&�d�D�W#���H�Q�g�d����"�d��������Ԗ&�3����X S�U��,�=��Dj7˗YSs�U11G�x����DfQ�sT�y�5諉�+��WZI͘�F	�+���S�㐑�Вħ��[U����Ӂ:Ő1�~���(��v�
���֗@��ѻd�V�.��o�y4����w��<&-��4���c�de�byiF?:�>�H�ʺ�O�30�?�D�,ri=z:�u���P��=oQ;oIJM�]�W>��"��G�f��B또6�H;�ٛ�ҙ�AT��RzciY���Kar�	g��A�4M^�$�-w���T}߀�AO�����\Z�G�<�\�QƂ��|8�)X �z	Uƛ��us���ۖY�N�5�^��X@e?�t�O�}�7Wu��y�+�L�U�<�udX+��u�Gs�-Jp��/[�-���F�:�C?6���M^UB����Q��O{L����o(옷��0��˥������=�(%�����D(@�̕��b�3��V}�W�������Git4�7���]�_��I�cH��7Q���ߍɡ��e�o����.Ld
h�V�Q�����8`��mY��c�}p"�ڕI�Sct �D+4OSɈ�⇭���6)>�ʒV�N�x�+O���z�ed�3�o��-e�?*3�T¹����Wp{��pg����|�q�J�G�V `sy�q�2� �~�-BV�g##I&yZ�G��3��Zug��se]\�F��E}����8 �����V�7F9�_�svt�` t�n��O�o��}t��[�Ӆ�z�M"�- [L)���>�G��i�&��јsv��g�mh[�"�������w*�n�M��
�,��p,xVd�QV�HU�����q����e[�Q��/�t�3T9���애��+����H2H�����sjv��a.����{�S\`�5��i�⃎�v�@l��?F���Z��נ鷷E��
t���j���I�źH#_joʤ���R����
x��F%�㢌`r��>I. D���F����i�O	�qj	�#�$K�*�u�.��w9���\7����9�k�ظ�+48ϰe�G�� D���BW#Zw�~ G4�����77�ri�5#�(0J4�E֚��p��aK�az�W-~�d��&ʥg��^����O���5B/ܴx1��������#A��{716��M-�`���X���+����t-���!����*c3�4�x��|W���,�+�% z������� ���lo:����S��J�7淴�2�/f���� �&�~�lz�M�݌]`�6�E��0|P�::B��_$p�Qxv`E�ٱX!�sO�?�/�jƏ̌K��J� ��愿ʫ)��ʿp�thm�R�
Ҍ?Q&-
�7�r�������P����Y^�Th��
x�&��� |th�!������G~�����7Z@�FFWx�����8��
�x,~Ccv�$�f��sqB,Dj8����$��R[-k��d�Z��em^0��f�͘��OBY��_���t��G{S�UV��e�yΰ��N��>�TǗ5�d��/Mƻ��+�:L�"�����,@��n��	����άw�0tD(�fUf�>��3N1X���x��Hc��R�f���#�����~��vȊ#6���`쇦&}�R�
E�$�ZVi�ushozi+�svYs$$������?Pd�XF���#b=�*\:�ָե{W�)�y?b��&�~1_aB4��f��-y��m�DOx<�ǳ��; 3��S���^ �Q��ڃRoe���g����(�CR*,�y���g��@�;��Ǉߑ���>U�f���D�&TK*�I���3F׬�� �K�t�"
�O�_]����/hؗ,�8X�/�N��Wj���˅0��{��p��o����Pl�呇�cxx�o��;�/����>G�D���EԼ����w�Y�7�Л'���[��v�LSP��z#�k\&�Ya�T�y#K,?Č���d�8�H��ve��-s8ķ�A'���4��äC�jTKW�b��,kC[�ҍ:x����Fpv�r��Xq���+ߩ*�c�X_�dO���齡wx]�2��� mZ����G�#��s��WdK��� #��o&i�Lz�u$*G�s�)�\'�-�m1(��<`�3o,��蜖вv�$��1腌�[��%#",-6LƢ)��;�Ga.�����L$�R���9�9�����5q��w37�*G��9��Iq�tr}e$�g�]���ԘmCm���A�g�;�6A�S_>j����n�,��Uن���ޡ��hA�}e #�!P	v��}L_$	� ��8���(-��M��:6�{��o�Д���0�Sw:�.-{��[&�����2ew��p�y��	0na(��*���/�#�����j8�<2$^�h�p. ���N���}�H���xˮ��9���n\8,x��*���+o���i����шw�uM��(��q޴J�et��z����%��I�iiqH0P�#���d�K4�TϥL�����Z��f�;&�Y��9���x�3���^�HU��v!��	�X��w}���a��f*���Y��=j[�S��xq�����ƥ���.2QڤW�[�f�؛�uL����[�ָJq��Ьf�h�~7�NR^���S�9ȣRJ�V�I�Z�9b�5ɴ�����6�'g��S�\�ȡ6q��c�`H�Eq��<�~�R��D�W��5��rw���W^��tI�$�7g	Y�� Jz7�	!-q�*'�'����Vg���# ���+�[2H�>�"\|>s�mh�C�br�?�"���h�U�����H@�����p�:�Del�� ��
.7�'=�1����k���&�bl7u���f-}�`l��-�ո�	4�,i�M�{ܑm�5J�`����jͧ�m��^�}���RXS!�Brc�nT�/?��pX���yC��/����mV���dB��GE��+6�L׈�g���L�Aȅ�{b��ܶ���sJ�n���_�5��R��e���cv�`�"�ә։cu�*	N�ڍW!�D��Ŷ)].>:C��K��8�� �g�c����%Dy@�6��BL����������	�馼����$��&*����֯b����)�@�u�w�c[.�I_N��c�U=lQ&̏K L!䳮'�{2�Vj�}f����B
$��R�c;�� �-v���a�S�g@�[Y�+��p��1��ŵ̯F9�+�����{E�eW�����+��V[�:��`$'�(������ĺ�c�*��4��J��~�m�h�yHjh �W�76K�梖ME.>�����Zs�h���(kg�����8GJԼ�Q�S?[��>^>*f3���/6"ع�OL�`������I�ĥ�%�RAC���8��2����ܔ~��0z"Q
	(ӗ&'i�X+8pv�)�t�D��(�4C����n�;=Ol
��N6�t�mi|���DՆ؛�%"��R���e�����TZ��=)�4�+#�T�.���A�9��:EIGR��{Fuqt�_��N>��=b�̞H��Sj�%�ﾆ�'&��]�l���*Cw���	z���,���[Hhr�ߊ�"�v�ّ��6�"zrr||��a8Ԃ�t��"@�l�0�C'm��Nu�gԋ���_%VT큮��V&c�4�*�M�$S�D��I��LV���`�oj���bS��zGF%)>~���:�	)?ߌW�|$�Կ*8�����Kŭ���0����C|ǡ�g�W"F%�]�?�K^Il��Y��C����m��/ӕ�T�+k�ˠ����.��9��.�K�j��,9A��|`?�t�&O~�,S�k�A�FX$KQ�=����q�׾{n�s�5|���m�突^B��B���6�AnH+Dr��̵�v�F��l���#��h���@G��^e�O��k����u���9Đ�/�ܺ5�[0�Hb
�J������~\*�GjIcM:kR��7~��5w���R�22Wz�5�(k����nm����ٶ�,*�^�����~� �|�O��X��I��15���-�&��{p�������TtD�X��aT�f���h	�?�WJ()晠	Q�*��b�Vէ��a��4+xӐ��;�a�%Ȕ`�j���MBN��{A	.����4.m���V�܆COs#�Y��/T�n��q�nL��%�,��׬c�O�q����=�&�{��@)��w=��&cຶBھNm|9�]���U�W~�f4��:O�`��v��n��h�僞?��clg'gl�w��)��Y�|�n���x�FX�$��nb���IR#-��2����zs
šp��|��/�D�u��(��9��R����ka��
���>�F��{�;��e�}`��?�_Hf(�j�sBj�7��$�hA�s �摀�(��?����r��朮!�6�1��;3�a�1��n�������,ܻ.�MgT5P�W(� ���8���~��SD
��)F-�\� 9^{L�%��Ng�t�ύG��z�i6?O��4�̚L�$pL���_���C�Q/�\4:��ei�X@��D�p��Ū:���R���<-F�;��]gQ� ���cl/$;��D.d�^�R��]t���j@.�R����`�|���v`��E��͐��<1<#�%��lSs�x��0��*�U�EI	'د������. /6�H t�{	�k�B�C�,6gb�H#ɱ�sչ��p1PF�Ps�ő{t��Ŏ�!&_�]m�F�j�LY,��t�����ݷ+�m,`V���oTL��86ϻ�<o6��'�C�"��o��]'p�(�fXT]"6oRG��U���q�Aʙ��:y-²��4����k�e*@���c����TX��7E�y� cA�%�i�[$+���n�:�����s���ֽ�����H�c�TS���s��������Y.���dk�-��Cx�F��,�!X	��Q�E����;Pnn���a���ոUJBg!��u\	��/N@�OPQ20�s#cŨ2���W�{�+P�	Y�����8�iw��%���P��_v�]��d��>2��?�N�~uo6�2��ן�Ql]�{�^��=m5��@�|I�Fh�1��I��zx�\��Ȝ-d@���9��ģ�u��슍��ǭ/�q����-8�D��q�5��al[X�B�Oa�C�eG���i���G[��%�!y-��<.�jQ��u�HIu�D�V(�����x�\5�a��TٸK��ޕp�~�>|��Ϯ9�?�@�ށ6�$����6�Dl�$��/���^tN$0�.���TX�����a��*���eX�}�e��>���߈B���򡴊����s�8�4x߳�/�,DCi�W!(�DN;|��ٛ����G1���1 �g��޵+s�3�Bj��nn^ =��H�s-^����}(�=��R���/Of�j�?!�\\0f�B���҅��j�F�����)�^�`Mó�d�!SOչ���$8� U��e�;'+Y�yڰ����P4[����β0�*��ȡU���@ڌ��Fi�S��1i�֛�T:����O������{�9��o0���Ҳ��T\LDk-��Ĩ��� �i��x�e�����9�����1�Q�۶�֞��P�j���5S��bL��:��x�V��u�:��:������-bPr$0�������b�V��#0r�����P����=ă�&�Ou3N�>v�d/�R�&��P+��l��]���}��vb��b"P�XNjT�Jh���Hզ�@lP!Փ���x�@�b^\� �=��߯�oѕ���3;�hb���o)"�,{aF5�F)��R�0WxW��G7��~���׻����J�{M�T��J0I���0�{Y|�Ѵ15&�4�	�nt�&oo��  X�p(=p����ݟ��vg���
��B�u��ju���Z��rh�&h�?�����M�`i�K��������x,��U��>R�j�j�3R&ڄ��@�~�a#�_x�$�r� G�8��H��s�	$�]t�wʉ_Y<��c��<��9���4a��L�t��Q��	%�ӝ��o;j�W��U�h�N�����Z9�^L���
�����4��bM�������`Ғ�
*��*]�@�[��E���
A1gOpٞ�	�έP��r0HN&��'֊M���]-F��a���U�wTM�g��"��I���Ll�������6���8�?^3�vo�-���w�	�Tl	(�9���|h)��4<H��3F}]/
m�@[���&6���>����WcE�QG_>�'��f�I�[��@���I��/�$��JVx�3���2~<�������V`>U�W�g#�Χ��A��W+��l��i�pzC�I�?��5(Ru4�k���Ψ�h��wK'
��V�$f��}�y��:S#Ps�0����¬�Zu,�������q'\�	]��K�[�>W�w��&����F����?���	�4�Fe1�(�vP\��F�uS�%����xH�U�p�i_+�T������mdpĵ���lQ����'��Y%�ʡ7�Sۿ�ldK��g 1����m�m�~Z.�`��M��A���{ 9���q�eʌ��
u��P��ay����G]ҡ9��V�XU�;z����6<�����Q�ⴟ�ٌ��w��{��+~�L&�:@����-��kQ��'�]^hj�Eyf��a�f�n���XTx�$��O�>F�F�3_�=�Y%�Q�^$STp��Bv�7��%$�>
�A��W�ũ����]i±��U�K��ALQi�d����U�h)e3U4��Qh|۠?u��亭�U5�*�[��m���iΔ�׉-:���GB�8�8:��z�ZT���N� �)3����Ւg��f������4[]_���&���bN�b������_�������a�����e|N��O�3���A��	�/b�2��*��T���p"�c@�a���.�8�u�w�z�f�V`���Σ\6Q���c��5�:�rG��c�'�g�κ�ɽ�F#OC��~���,��	�Y��*ULO�n��{aL�G�?���L�E�>+�y�)���	�k7���1�!��uѓ��E#=����0�� 9<�V���1�~���'}�|��&�T������I4s�*J����U������Gm�����7XU��F��(� ����F�K�BĘ��<�ЗN����h������N�/��I4w6�5slF�wQ}��:c/�sh�W�8ߒ$�v'\�qa-��!���Փ������`��Bw�����}�d��b�kVcZBr�5y�P;�}�	m?D�Ui��Yt�~>�k��|����x�;@�a�i�h	�Gs�$&�K�oU^e)c;@���UwwXn^�v�$���@!m[��qϋ��E��F4���ܓ���uQ��[�Q�u�CT2r]�e�s��*�~�ƨ���'>�pb'z_�����F�S=t��J`�AT�,��~L���*j)V��S�?��F�����JuLr�mm��G���A�L��v��ܼ�DOk��6�U	,��v&�V[ �B�3�ŉ����"��ѐ��m��,��Ȑ`�)P�b�Ey2Z����gTܠ`�
)��7ף�t/�
��b-��I��Wci�YnӤ��L߷���Y,�wxȂ�)d�M��%��+�>WJ�^�
��V���^��[��-(k�
y��P46�{0�F��Uo]�w,\�t�&�N���օ�B:��oe�����:p*�#��uN`�-Q���u`��K<e��^ٶr��ܱ�θ���Q!��ĸ�� '�@K@�bNF7%�ߐ�2-�U��4�W�޹�q �Ώ](&����t�܊=/+�v�3#( �Z�#�F��lKo!V=�@�I���l��6���vf�&���)S3٭�P� :�����R����3Y�߷`�/�AF����R#�gO�jr]��c���(0l�jl�z'``}�d!��1cw��hx����.!N�8�OPvOk3�a���+-�P~�F�8p"������>���<6�.��µodX��z]A�!m�Z�qX�H0W�_�FW�4�X�������|6.���rk9h������G��f�HF��H3q0��Q��J�16���]"�Ϩ\�,����$�>�V6q.U�^"x��wjlOC����`P��%���a?Z��d�k�+�b�kB	S:��|e[M�MCr�!�Xr��i���č�t)"��db��HK	�;�o`r���!��{�8���^��k�yxw��W&>�uB	�W=�����`ɻݕ���o0ל�g��O!Z��nd�ٔ�������ec^,��l*�Z`eS2���u����ygĲj&6Ed�/Tm6�S�;i�n`���X��)��D��c�v���c�{k��}x5��j\�>i��L@W\q����o9
K�P0�?�/h����2��#�r��+��孶��&*�����ts��7�D4omoX�O+������c?��.B���EMSY뭘��h�� ��]�pT8�����˘ؓTlz ؛+�k,e�h�g������-�b���_J#�$-�h�ѕ���_��W�i���XQ�?�HG���9Z溄]�ȩ���_%	45�v����kf��:�s֒��T��h<h����CE�hF�E���;$�*���[�Z�Q��b����R;ٽV�؝�)�u}�,��4���\���
��~~zm&��@��p�tˈ'�mfni�9%���u��)�}�<�	qp���Q�ܲ�M'���;�I�(�[cBqy����L�>ڲ���T7S	�dEo�.�_1��kD��#zj�G�1�q�.��������x(8ã}�۽,�����sD�"UA7(�[�(`A�4�,ը�!�AT�E(��tjr���R�]V��m�^��qjX$�-pm~��������V�Ÿ�vX�q�/�xT�������z=_l���"Vdյ��)�H!*OHt�'_��R�!�R<��4
�#5�����Fyd��!�F���k����Y���h$K�wY���͏�f���S�����%�'�����|ud(�W�[�`���5e��/~g��SV��7am���p�r�3y
�;>2\p� D��a�r�`n���9�V�g}L3���Z��6_B��p�2���!+���q2�����|�I~�`���n��y@�(��J���>/7�d��+��˻ ��'�ѷK�%���cOl�c��J���n�E,����z����q�A��p�W�����Ŭ����g�D`����C�U�hSCo�+���U��ޅ¼��UI,�4�NF<�7[ ak�b��$~T�'�������(h���eeF���`�������h ����Y6W^D�r���H�_����>B��G?*����o�T����`O�[4:9̝�b}�OA��w����
�*�٤�}-]��d<U)N�Ve�6s>)s�ʮ�a\�7�D���|q�ݓ%O޳=@
�QYt'ӆ0�E}�
ΩsP���*xnw�R?�jˣn��[s�oe2w�Q&�i��`T�no�L�Y~'~�G�U�W�=xl�侫�ךxG����d�,�4��,���'�־PX�T���W���<o|z���d��0�i��3I���EI1ye���O^�D����G��-�{�¼j����:#�g:58꿕7�Wh��!�nH�sP�Z�q�E��`XOkXт���1����'���X6�IY-�L�0�M�|46�SW��3Pr���]�8�zX>ߔ�h�>{*4" [�!�j]���s#6���Ά­����RQ�`���������rh*F�'�,�̣|c�=�,��vW���q�T�kL*+�G�G�y��`�E��@FvZx�4��N�a�k�Q���i"�DK�h�����I0� 8|㊖*`o��ÂAWBuu�~S�H�rPL�{GA����B��m�9f�v�{9�S%5X.�l���+��@'����o-D� �p>����X���
��v-��^����>���i����&�,�I/��g$�>�V��I�I0G
��	s!F���� �Փ����K��SJK\=�fy%��oz�2�X��_��O�t�S�{:�}�q�+����Х���s>�@�%���C���1�ѥ�� H��d]��=9�[�(�\X����)�i���ȭ\�m��H.�3��
ptJu[ֹ�u�D.��UP�;�@�U�|��R�ѹ:D���h�O��!Z�_Q��#.�_���å��7T��{���{�9��*��/+�^irQ�VNR�����X~t�˷��37v�0M,wJ̛���w,���dʹR����ԓ[Ѝ�7Ng��9!��*Ӊ�28�F�G�����f�X��n�σ࣓��\Hd�D��+{(`�B�!� 	�P,���mbΦ*!�^d�[0�e?���J�PU�gQ(�k�3�S���L8���vmq+
[@W牚�.�اk��}�q�
�o�j	"��Cx{#��QL�Ҥ�����g�\k����w����X,�K�LFm-��I��ֵ����h���!�%y�'��YM�&��b�u�޶��Y�K.��)Kn�`������|�8X��
��M F�I�槆�������F�{���9MV��`�3�]X����b�QW`��j��%�u���H��rs�P���L����:��y���.�o��l���Tn=�u��ݑM�4e�Wn���OC�3ji	�Zm�ld���<� �A��ؕhe�z���4����� QK�s���ˉM�BP�%�f�ǣ������V��o����y$�k\h���Ҭ�F���Z��c�F<ڽ7L�PT���\9���G��z�S��O�{�@�C--�s��9P#a��\Q~X��$8�(��4�$,֨���Tɜ;F4/�(X�i�0�υW\$��RY�(�(�
cbp�( �:�agU��?��Fy���#n�i������Xxx��1{��R[��jo����9���.��Yj�q�A�eM|�\�8�J�y�_�>~���I �lz��N��N\N�Y�`��-�EֶH�.w�%M.��	&�����3���@`��1 �Wap�����e+=o���^_C�QUJ�Ltlt2�O����W��Rv��<*��~P.�9��=���Qw�{�?%�ݙ�Δ�(�r�Da���4U��w�5!��CVy�eA��2�3�����}r��{g%���f�m�o�X�)�f~v���ʸX��dT�e����v�_0�k��}��˿l&?OSf��uƾ~�X��km�����v��9>�K3lp�ٙ7� ��q�c���c���<�',��a���D}�w��x�!�r��E����r��?�����+T4��?9��֡�,��e����F�|�Ӹ��ȕ�����<�Ԉ��R{��*v�Qc��)��gS��
���63z"�Ԃ���[dt�*�����K߳y�yȹ��[�E�� I>��U��U����1�G��N�B���ԓ�
��.�՝|�D�(y��s��Q��,`���)F���9�H����_�E��; -e�O]��P3��Ϣh$�W�bV�t�`��h^
U�mr
�PqȜm�����)ԡ��)��'�CA�M[ᄎza2���jm�6��8d0��,{R'|�z.��S�>�!4*�vl`����	+�],���Jlne����M8V����U
�30������P����4�1*�lh�{�(@��?.��� �u�-�(@O(%GB��U"�E��X� �}�+����7��+�Db�L��Oٕ6/�.��)��N��u��H`����@��i^�4hkC��[����u�[�MO
�Xv���,r��e�|�(��!8�BtN�\'��T	��'*>�Ν��pV�w&��5˃e�4fjp�u{�ć���ٶ����d��Tԉ�,Q��\qUH���*P�D'<�Gw���"LTO�'}�~�p�R�3P��0"�oY����0�Ѕϒd�)���mצ�ʑJ��g�+�Ô7+_/�|u�\_�� �:�3�y�h�(�E�GB���g�����L�Z������m⋹B�ޡ����,��
�#z=^��M��U�yvz�-kS���e:%�a��r����4��`��N�4��JȪ�!��uq�ve�@ܕ[�� �:����DM��}����e��+Ȏ�my��	�� ��C .��PA�F����"���s������~}��,�?��*]6?S!�Uj{�PI���nC`�X����~/k*���X���ơ���e8V���N��oy�Y'��1FV�X���)Ph� j���o�`�I�kU�l��Թ6 �Ǹ�-�m���vd�0^��2lmpyt���/3��[�S �7U��c��;NZ)���m2�W�A�y�ҩJ^����`��J����ؾ�>~�;��^�:�
�|�Ƒ�F��ˇ��bcԐ�$'gX�����Avl��S�S����SU�X{.�f���)H�� ����-oD����@űn����c:#l� 4����ۡ���QO���f�u�?Wi�|��*��������
C��8
0�(�L��q'��z��ڐ��]������;sW�Qz��!uر}o��7�����ab"���u���w���_]-U+PG'�$8�d���?�x4�3��9�\�ʂ���5o�f��:I��J����˂akVLN��.+^�V��h���c�"騌)�d�kr�NKd"c�-�t��:o	k3T��	Txi;�M�z��B�x��:Ήp�3)�rXn��2C�v��>�Y"��{��[-c�
b�^zh�%���u�~xw��2��r��H#�y¼Tf�"GXH��b�^*_�GX]��VW_�~�%��
yB���y��#�!��̶n�c��[�#�}B]�+�b�S�#j)6���R����Z�E��6��W���H���#ͧf���u(v�Ԝ�O���߱z���D?C~��[4}Ir�lz�����H��L��b4�3���j|L0C3�$!{:9g��3�����NAnԳ�r�1�  7���9(����MYT��9z`�4�e��H2�ЃHc �۞�]޿n�$#�r�������x�W��@Q�fY�ʛ,�p/,�y�}02��G�:O/�&]�?�)(X럴�m��t��q��	j1��p^9��#�d����/�W��:0v�C}2E��?���q��%0dȦ߃7���1�aO2�F*���}��Vn�7���Ջ���� _�����e�v�'l��-4�%m�H�������W��gH9ݲu�A�䰳�$��?N�i��4Jz��F����dl��!�C78� ��R$*���Oغ�/)��|
Sy]ɲ���E H�
��L��L8j�K<��_��#�y	�(�V���t�:q���/�9�ՌT%���O���!��D%+:��j�54�$z�i8{j%q��X��Lz��_'���1�����%�»�CE���/��![�HP�KpDg��q`���N�����]��0uG����3���ƚo���T��qX��5����weRA1���P����1�}�,m#���^l*oa^�xy>׾GֱL�}��I�/�w\�~IA(��;��Ե]ZJJ��\��)���cR���@�-Y�W�K�ӊ���LL���#�ف�%8cwP�����|V�`���&f�3	�b	I�K��LL��ȗ�"8ݽ�?R�Xʈ9}����j�|є��eu;�r���y�([6���4~G�xIs�2���Yq���������{�3�9�Gs�z�!N���t�ޢ�D-�Ww����:V-EL(���'����gE��:W%��-'�[_ȁ:x�տ.=K�ZOM6�JQ�_xE�0ㄪ0�s�$�=�G�^>�
;g�e5W�<۝�U�eI��V��&\Qm���eU��3��`��*�t���s��p����x��.E��.���U�J#����e����Rrd�|�$b�4��[�]b�;�`�G@�~���ȋZ lI�RÙ$�2$tp&5���uo�\�#��w[N���D�d>R�d�wVk�����䯠K����[�&���x�����<~�;�����"�1YM�u��T�����	ў'�*|J�����P��pH����op�$�����s0O���F��Xw,7D����V�!Y�xI<n
���LC��>u�U��ق�UW�̝��wErE���#;%��n��)�Xl�6_iσ{/,M�zz*AI�59B�h��=d�
�o��&Ȑ�����R2���T�g��E׃��N�c�)��� ��p�m68�;@���Bd_��e:V)���W�?�y��1&)�3�1�D'��%�h��1A2�PVՇ06�Zk����Ʈ%Ht�{d.��B�����(��?ܮ>]�JeM��o���-\J+���,����"0"'���'k���nz�֙v�Sd����
C�>5�݀j�kO�Z���z�\�ʻ��չ����$�	�	h���ƭϏ��/��İ�r�+�3z��Q�Y�S���(�����>FJ1z��{�[ܙ!3��׃����A	��q�a���ъ��0��
ޙ�F�����Ϲ9��?	� �'�P����M�f��<�H�^&^7P��M$�v�I~.����3Մ�m �X%v,�\���]�=q�W�m�t8᪠K^D	|�s������>7���]|_�=�ܣ8xV���c��|Y�dz�U=ou�1�6��ՐXS�;�/�z90ɿJdiN���oYWȺ��<K6A�-�A��{�k(�c�Y�ǉ���G�}��6?ѲH�-;���0�c�#`3��`hQ�0�g��\W�	�DLg����ѠJ����O��#Y@u������`��x��ք)2T��`�H�x����9(�HZ
�>X�</⧧�Mch�}<w1���&�kC��J�O.@�A̐������Fo�eJ�#��Ƞ)|ȇ̑l?�3#i��}�k��|�iR�3'��f����ZPL��/��|=<Y�6��ÊΏ�(B������p��W$�$Z��wҸW�5�	D]�ԩ�$� ��vTRY��4��+؇|-<�㾹�)����i�H�宋�X+��鮿Y�%���j�VJ�Q˗L�I��ZU��ץ\�B0%���6������&��kL+�0���+�=;�};l��GG%5���ʧ%P��p�{�t�߶o��j������ �G�ǆ���d������Kj�{������sf�����fiC��J�C���Eͺ,��_l!�nm��jA���tOwO�F4�������Vys	ƒDˑ�����`GƧ��4�ѲF��#
����4���j�ڂs��{a�[�C��/,���)_.��_�ʧ���s/�vF��巜8���X0�N��3�h�9&�����P�i�$�ũ�a��!������J+"����f�S�Ji�ި��N~�_���)��COVH���	p�.�6��nr��,���I�T�=|������B�Y��`@i�>�P�"��k�1})�Vz)@��w�'���5�Y�jn���6��"�\`T�]\։o��-&������>�X�n�������4˅�ҋ;sT�S=�$0Eת΁X;R��==�Ӳ�������w���&c"�rt*/�'�7��O���7��$=V��[ȡB�������t䨘�j4��7.0R��萪?j6�e�bg��i�8#=�I���9�v	]��aBз����G���}�C�o��` L6/Ǔ[Ĉ��t&܏V���A\�.>S�T3$�ڰ��=����30���f��t��&ߪ$Q�E���/@*��p�`l�T�i|�(�kI s��ϡB����B��)$�l���ZAn�S��0}DC|u M�H�_8�U	j��mJ��]���hbF���4�z��2� �l�O�}��	�
�����2��B?��Sq��쓅���9�<��q52CBk �Yw�Ng��"�f�c�,�z)ʾ��L��;Ƚ0�V�8�7�:ͤ���!S���lZ'��]�I7'��`u4�3i�K���c�Ba�����·�߯�7��_Ө��+�,9z��QT��||8��k�M�E�G^�
��I���cnN��S�V[�f���1[��Y�-��<+��X��a��-U�vݦ���c8X��~�ߘ�x�p$nǷ�\��� ���C|��R���3���w�)KN �n�έ\�<RO��bn�7�a�C��`E���s�n�xϱ~���w��F�����Z��ƧG��~?g(�,5t}Cx� {����`���ĭ�H�P�:�"`����8�3�?�˲�7k$'ZQDA-�i��L��ΈW齯cx�b��JL�/+��G@l�œ(�"A?�&5a�^\���%z�~��<,g�^�6�K���p�_��]M���O<qGZ�hk�%�,8�*SlMQr�8SW%�-)�e������>�+v')��s��Z&��]���G�߁7���J��&�֑�p݃�몺���� XD����c涾�ca����t̆9Q���И���6*~��ȓ�Z�7���k_��#;���`�؊=d���J�O�Yl!��oa���x�'��&��-5"�q��L�nOSS�檨��V`�/�#H\�i�A���`c��$$�g~ڡ�w{(+&fqh�
�]Ō��qCê?�_bs��g�jCCT3�Z(����ý~�X�-����0�&"׽Rg�ݠ��h�����([�9�Ĩ��4_���X����4��:�0�i��x߫~�%�4���ҧ4R��r�Y�<( ����omz�a���׀��X�^�6�CX�˟� ���:��N��_��Ս���ިiXf�9M4��-�p}<{ ��n^���-i�H��E��I�x���y#� 4�zG�s�o�ڃe�` ����0��{�)H�02^���UI�^��ƹ�zO�H�FA~Ac��*_��@>
�<���l��d��2
�pFB��6����I�u�w򶂁�m�S��wgS7��(�G$-�U�BZ�C�F�o�Xa}^��$Y�4	�?�J�Z�N�gY�]]��]ִB(����,H$����\p���[:�V��4��`������[h�g�J݀wo������R�ޫ�	��>�іDqt%�G���b:��>)��5L#���J�~���ږ�,b};���/����"�((=��e3�����֘Ae�&,��{NB*�p�FX
��H8ܢ�KL�4Ϲx�СzC�p@ԅA�T��UK��金�Me�YX +T ���\�uu�����m�	�>-k��/^�����5��Q��qeσ���ko�T�L�U�! �f);k����+��������5�9{2N��r����4It^�|�+��x�t��D�����*������� w.�!X�����W� n��B�Ry�El�#O��͏�
[��5��(B��+\s�5�}45O�,���϶l�y�">}(^i�<M�У[S�U�9�Q���L�l��/�5�����MK��rA�R�9_EC"v����3_] �v�Gj�&l8��;yi��� �@m�޽"�Ԓ���և�%}-{A$X�m%٪S
���[�!��t�w�J�s dqT��@s�s8�r|,�i ��Y�qS�:F;$5�6���#��Ie �T�!)<H�Ao�������,�����r�t'b��z�BWk���W+{�2
�����ԈR�'&������C�bȥ9�T�	�Ҝ(&2"�_=�L�I��W�d�9J�p=���a��ª�8�"	�]+c����\��CV4��I�{�}�NM�ߥ),լ$�ˠ�B)Ǥx���Ӿ��9v��k�3to���8��2m}��&�9�FL�PđZ��y��|��3�@��N��{C��`׽%ԅ9YV�n{����Nz�@����dג81���2�Ӭ��y�H1P����E�Cu*��<;�ܦsn��*P��n1$��% ����3Z��A�Ҳ����e���^Fj�'�è����=U-��(I�*t`��:ع��͂�$��W�J�2��Y���i��ȵ�ʹ��Ҧ؟e�]�:иjK��?�4� A���I�����
2�5-hO�=�nN�Q�/�y�_�c�V^�z�J���!�� 8֖-	�#�&F�W���oA@�Jï���\9l����e�VUT%,x~���:@!f
�
���nf�I�l��LPF��T3pSC�ByΠ#��nk����5xa�l���N�l~���`�t�F���Ԡ�=�P�I:���䋸��-���(���!�9�Zy��)�)z�w�4-���ׂ�q�y��R����6������
�h�@ GG�������0@vY�S��M�R�R����L-����I�/��X���wG���zg4��<g�r��!�Bk��uK@Hp	����"x{�qߵH�^̳?c��(ܨ�h�Jm�0\�N�9}��3E�v±��O(6���s�Q�����jcn9^X����	aP�x�Qj��
�ߵS��4',��t�Is]��Ӻ`�󚏟B�M�^]����
#lE���t�ҹ�x����e��׾���x���@�������G_��C+H|P�00�|r��qb�,�y|t7|"UM@�!_`c�H�q`%�>2��� � ����{�$Z�i/)#Qp_4��B(�^�̅
-�1֥̄A�m��N��v׿+v�x�բ�"�7
��-�S������#�CLKb�>L��Í�x�#���z��|iN�*��zD����Ic]�ft�A�p�􃚋���K���d�@���.1�*�9KT���U�N��T�g7ô�RwS�pH��:�F�4��׭���>H���BFk3�h2�i?}J�msr.j�EWJ=�==�7�H�����_��8��D`��
:�S�"�:���s�LCw����Q=�HIt��`0�o��JT���~~�f5iv�S�T�.�C)�E-NJN����P��]��,j�cvB�l����{7�	{7K�tU�@�{�	�2h�1j)�;Hb�p�(�0�����.��i>�-�9� �j>�Rg��c�iG�L������9�3�2��ע�e(����+{>¸�Ds�}�f�As�B^󮖘���Q�ѥ�C�2�����YM�T}II",lF���a���80㲀�b<0�ڛ�<b&A:
��/�ծ�R6�7�L�JM�=�[�d0��3����.{�^������@��W��,���;�*IA����x8`��11��g�>� `����p"�l|���µ����7{��'�o�q��W��\DL�^^�z�Ý_�D޺j6t��v#.�.��@�i�Eè٘�?ɔBƼ_z��
�U�j�kC9��Nߞ����$ri�jkU4�bo�v^��EZiC��N���e��+����מ�V�r�5��w���з��j��?ׯ�8�{:!�N��F3���k����;��a|��tЅ;�9�ܫ�D�<nr���e9�d���y�W��x�g��B|<���θ0r�=0!e�i�#�k�;&��&@��3�kk�U�II�f5�	Odz��l��m� �L)�=9dd�K�K��UD�(=�
nb0����#Da�TZ҆��ha����M��_�G1�KU͂e�R��RX������.��
�hhɛ{�~�e�x���!͉���b���d����Zq
�B��jz��3<�j�l�Q���GJb�v��i�t�����(�T��#�<a�2ґI���,k�8�a �Q&;jݔѹeىs"1�d>Z���V��lS�޷��?��-�iw�"fc�_$u-��V��RhU!O�/T]Q ����>��K�=� �L|�7�("*�wj+������EC�M��-��qF3۵�����s@H�q�O��TL~�5k��`I��ғ�K��PE&�f�3Xl��v���,�۷��`�?6b���ӵѾ�Bl %C����!px��iz�	x���--6Aֶ¹:�py����Aa8:�5���:�I%�P��.�7�[�!d�V��Pn���tvN��L�^L�IB�Ҹ��n����8I��"�	�J:����FՑ�+w�&N���#h�kf�~�GY��X{o��"6�0D<}�f�	����W%i���l�ʛ\�k����9�N.�oS���}RA��q|B�0���~i~�0>���Kgݣ�S��%cr���ݲ^�����2��	"��j:�'ׄ�)C-�5�!� �K�����K���K�Ч\�hb�z�0g�����X/u���@����Y<<R�� d6��w}�2]�T����<���ņ�P�7T3Ym�����Cp�e{��V��?�5�l	�l;��9D��#6����f�ъ��7���Vc�_Ǡ�P�g��	Ͳǲ�xҡ�s�o�<�=�:��ѣ�9�ল�z
�߽����;h��E�̍���A���xs��w�ŝ�}���wtn�r���!%�S%I6�3eI%�����LL�IS�k�=�%��5H�,F�Tt�H���?���V�ӚW��e*ʹ��+���������'w#�ZQ�U*�&ȵ����N�]E}�se[����4"������'�M"ZXU����I�бT,|��eh�+"�b�����ϝ��z�EiN�%��l�	�0������=�eƺ�j8�bG16ۑ�B�ܕu�o>�+��3ܐ�j�6����\��$鞳�sfC�BT�GؿHWO|�9���S�b�2�@Ǯm��K�c�\N�TH���PUL_�=�E�&�[Z�泊N���vc�5�;�y}�vr�i�<��g�ř�"�^�f���)Tj��T�L��g�nG���A�;��!�U����E�B#Q˃�*J2��V�v��k����u�/�:=L���<�������r��-��;¾L&��	�^�@�z�=�͛8ԭ��u7���9���|+�@��5v�G���&V�s��(nǶl�()��|�7\+*}�hǣ�UD��QH��v��
�P�e0��S���g���[&c$NJy���\f���s\�.n��V�`vlOlR�|_3�[b��$y$T�Ab��*�� }x_��S�a��h��h�=y�x()�}������v1'ߵ�9�o��%�~' T���K��%�Ds�3�b"���������U�)=�f��:��Ϩ��x"x�L��E��}��@sPL��W&|�l۾�)k��������LO��D���ɫV������D�D���*�E�h��r�C����m"�FO_S7�^��u��%#k�0!�& ���O����-��/h�a3����M��N��|�ê$���ܥ�� � � ��z�o��g�"��/��y��d����e4�F�s���8L�����)���o�Y�f��|둎�N�=D� �nD���f�|��l����&��9biJ=~3]�b�<ۯ��1Xݐ%/I3|��N�����tL�H�Ǫ|�'<���$_J�P���=q'3�Fm,j��M:����e,�(�}�a���xo#�ba����#iisY� [YV�чK(Z�s!�fQ����ۈ]&�����)�sJ��:Ě��U)<�Z�״���x�-��j�Ƃ��S�{� ����6���S�[@F��[Ӄtz"�ȅ���{�m���κ�pN=7�\��Ɣ��ɼZL���f���J���(�w�ɟX�2_%�e䤔D~y�٢�z~�W�.J ����%��B(�J�3�@�B���������4&���2܈��V���I�R�>�G�E�q�j��� ��>0�Kx �A�)��ޡ>���������V���DZ�d.�gF�������P�3��ý�	L�_~n��a��������n��p�?H��s%�������z�B�׸�&LX�:>�`Hp��v��J���e�^c�=���do�̺]����h:ӳi��"�y���.针BNE�I�}=��-~���YޅqJ;��<`�ϸ� ,���8��G��=��z9-!f����E�T�!��ᯍ�&TE.b ;r���
�n���\7���2�q�-ڞ��X��1��D����}�5�ڡr�K<U��V+��O2��9�0���{�(���)H��ҍ�O��e �\rp3��V��Ϸ߇"��P*�V���<�,*��l� `Z�J�O�]��\��sg"�����79G.2H.U*�a�'{П5HYl����9�!<�W��ku�W1Ϗ��>�v��ܗfݍ|�V�t���%�2�n����J2�[-��#�W;01���BgA[s_1Rs�ĥ��}�SwfL�hٞ�����&����TJ Ê0W	7Un*�1N���4L��Y̆J����?����w��i�>�bp(w-d<^z���Y��eD�����ُ��q><L��s����>�����0a�4
�ng�~�	��)>m��bkfmވ�ys��{���f��m�@46��І�nm�BX.3��k'_2�Tr9��H�������7��Ư�����7�a�
4���7�Դ�z�w��A�������P9BWɦ/���t%���~Qi���+�n��U��o�c�p]E�"��}�C��!}8q��XzO�
E���|)<7	.R>j�^� [��#<��rdzq����J����]��w��q�w^i�'%��R�
�������3{����A��ؓ,*./E~�x��p�#��gW��ƹ��)/0��9J0�������D��(��pM��;����,�R�t� �3���:.2T�ۼ�ҟT�A��"(�yiov�p�-1+[vp�<]y6D(a���pӋ�y�5Pٜw���8v��#3�ʛ����L!�F����m8��.�G�^'�ZX���$Gd�w,?�N����@$g�<,�����k��h�K��1$_k�U]���-����:���g+����ϥ���(7;��R}�:M�p�bV�ՊUp�7�@3�۸ľ��F���i��9^������G�Qʒ�����6����6C�Ǔ7�.X}K���;�����oF(�uQ��j�D� �~pfCA����U��w%�����5x�����rʻO�EE�3} x�0���5P�
j��ݼ;��'��g����F>���ͬC���A��z�����-K܇U��_�CFp�lǂ�u��Yy� #+Y�h�3��aj��f����ӽ��sb5����k�)���ܳ��-�G����e?{U��c_��FV��
.�z1΍�!x�:4F��Q�[dgMP��cL�o+����Hn��"�kCFS�N�@�7���V(�,O�t-�\af^!w�j�{�y����'���V�����N�{���[FM��2�D�0�v�~E�ӻ#��.��t�`�w�i����W�֒�C�	�u�<���q{4!��m�s�ɂ��
����3K*�F���(�������lU!R�i��'5:q�F�TͪA��,l�|���*{6���?����р�9��q9n"���_Ʌ���7�5�,e�SSe�����񺶫�\ݒ��&�GF��=z��+Ր@��4���ꢚ.�����	�4'A�AKk�b;e����\��\����?���h	^�~1SX�&�� ]���1��Ht����U�w�C��,���yy�Ʌ ��-��J���C�L�%u�Й5p^v��L�21�
�B�K�O�G$�����t�_�B[�V �L��o�;��i<Eﮪ2v���Yb�${��,$���M J��dXGV����7���`̟��wk/k~�L@e��!�<A^��Y���K0Y+��l�R+�
��s�d�3��]Xp���'��j��n�8�T�z�j����i���M�\�r������w`(&x������L6V�,�l[���b��~��.~
���	
�hj��� �D�C?��(Bc�\��{�Mצ�¼C*&eV��ZO�K��c#g�+z31z���.!#�`c,J� X�ն����g���6`�c���)�����T)O\�$L���n�l]^ձ	3o��] �LS�/s���$Q��e��r�xx��z�g�1^��)��
5��jf(o�{���W�|�j+�2U��{%g���$\�ktQѶH՗���1����J`Y	�.]C���VLZ`�`Y���ׇ��?��j�j��v����fd���Ż;�%oȼ�B����G�`��Κ�A����=� `�=�s�����!�gJv��,��ni��������A��B���*_k�4d�i���%԰�r{�5G'@d�/YӐ�$5x��Y�V�x�.��6E��ہ��܊���0�'
��� ���F@<߃q��%F3ٺ��U/�w������lɲYˇ� �*�}�nyE����A����8�6w� J���ԪԂ
�2Զ�}�fխT�ڳ@`�Op�@��:���Tj#ݶ esU���Gk��	N�D�A����L���8%���x� ��bJ�ώ��lzLI���;��b�U��H���Ncs�=�������$�ZE��X���r�  G�*�#l�?!u��T�U3K^1�-����,ׂ'��:�x<%�B�H�Ǟ���e
iM�����sjM�z�:��q��M�|�Z%hη�+����_�h�֍��|��\�e-�����^a*aS��Y���I-�F�����tt� ������n�=br$���MX�)���Q�4�������;��Ϫ!`C�,����w��<�8�������4��Î�(��6�����O7� Dj���@��Xl�����h^;��
U�׈���=�Z$;�qgr��C��}�N�m'U��y��b��f�%q�0�d^f#U�k���� �l�~�����=r�"/��_���5Ӷ�T�J�C[���?�ԉ{�.��򁞮s2ɩ�Aa�5��r՝�0;��S��ʀ^9k
���xloh�3M�*0s�Z}�{�X<:Gf܃W�J\�u�u&�9�Qt,#Ǆ�=�tq�ѷ�cXծ�p7�`�CZlLL�9�zx/
��χU
�<�,
������s[�)2S� B�(�Rxz�ӷt�-2��B���[Բ�B� G�0��NE��V%�p�E�]�h]�uv�/MW&�>��\�i�D$�l�������!�~�C��:�w�$����L.�����eCb��������[��+im!W[�:t��lt;�aA(�����D�`�,d��?M��.�+���]��2ݐ��p�2TY��U�r���>�Q���D���&�6��%���J���ec�ͳ{�ˁHO����UM����Q�0��G"=�T_���
3�N}��1�LH����a;c������i���4WϹ�Vc�>�W!�F���Ǌ��D�Vμgb��k�Qn��{��)��%�o=<����ne�i̴�]{b
X�_��������O����i.��y�!�#1��	Z�;ʑ�>+�[��1�(��@g�NE���N�h�<7Z��7Y:zY&�ތ���be��Q��"�F�<s��C׏�`=��#��L��_��X��k���#�Ȟ�c�3<�5dDN?ͅ�p%��.���7��X�f��y/O̪{�{�0ssJբ�f�A�#.X�N�|q�Ĳ�a�4�9I�,�ʰ��	SŇ�����ߗ���fr� ��y�F�"1��^��T��a�\]���Ք�
���3�y��<���Ѽ����8�0,���"�O\��H�\�I+:������y.`���ۅ�K�޽ۗ��@R��������z̄9n��
y��/���t���U$��4�P��R~�1n��v��zo���U���E���T���z�Mc�������]d!m� ����80��G��풴jQ�Y;i��E\�bzܞ��O﯏̗K���4O���Z|���׉�,���|w'�BC�h�n��&���}w\��@�l���y-�%�ƶn�����S���*��=��:o8�u�Y�X7�� JF���Qr��Y�#��Ne�TK�ޠ�cuL���6J�G��.���������'������V���逤��\�dF�\	���e�ň�5�����9:��"�tD?�1V�%�$3qD���N�B���u�[��I�X5YQO�u\R=�ӡ�
�8lb1���+��Z��"��W�)���|p���j�B��pt!9?���ﾏ"VP�U�'b�Q��|����j�����\���74f%;@� <�ʅE�:�W돓�]��!���;zc�I�>����!������5���q�);���#��q�H�;�}��Yo[ZQ�E�5�'S��Q?�ҾN����t^2ϧK�ɄUw���+���#;�b��`�n�Bpl�
��{�BY(�\�	<��|�+�fw���׉8���p#���j�^D;�~	M?J{���ym�s�|(Mg!M��8y� 3�h���'����	���f�:�(�N��`��^��C�2���B�����C_A�g9��vq@�l����B2��g� ��x�2��/�#��C�S����]�/.�9�jxX�þy�6m��q�-�g�*hRC�&_���ɘ�_�:J��C��;.8���	���<DE�sο�»b�$��V��x��ф]��y���5'M����O��F�q7;`��ę�"�p�H(��jr�hl��G��ՠ�Q��TF�Y�_<��u�`Ej]H����+|��ݝ���[�x�?�:��l�1�
�8�cu�%vF@�N?.�d�h�{Ļ9Ԗ��p��f�(ԉt@	��S��[��ɲ���r�M����Թ�vz�
Hϴ�]g���Ϭ�����Y�!Aҥ����`�u�)�d&�nP�>dPC�NO����9���H7�'�P�g���
����/�a�?��5������|�l��p�⢨�?�v˵�>_rE���HؑO7 H��8�l�ʆ���)&w��<�{��1`�%�9;�n�쒟�/�[�-�2��g��$�����zOͦ��vu%�s��O��u:�/���\����Ԥ����޺06~8tНc�,�ϓۦp���WA��(�M����nJR��(1S���P)���lŚl���,g0O�+�i�x'��"m��MTi�����qܮ8�+V�S�E��6�fk?��z�����g��@T`����T��4���P䕑��3�U[Q |X�l>�p�j{\lͳt�y\[�e^����H�I�?}��?�����C=��%�{���S�9r����/����o�[()�ᑺ�� s����*��-f�����6��\�1�eT�N��
Wp�X�~�|���m�d��J��ȁC��(v�hӛ,<�/��ɷ�����L��x	�]����gd��[�P�o�����1���p��bQ�*�����ӷA�"��G�/Ā��D�X�ev��;�3����<r��ځ)�Ў��n�4��4@>⅌x��|���#�����f�ӋuQ���f�OmT�C��)�% tF��m�^&�?�ϡ�z�����3�|Y��nk4 ?jXI��PUJ��ɐ�2B:+g�6D^��HS��/8\��!���Yҗ��Z�q�R$ �Ji�������M(��8�k
0��T="Xx��E������m�6�۠��8y��������0���3#�����b��#�� &���[yz��J]�аW�=��	q�O"Ԣ�O�,"4���~@j�ap��ۃ_㲎b�r�Ah\Y���52
��[�6��&*���;�ᖮ��2�L%a�j���ve	�d�C�y� +���FE�=��(o��3���@7��{�D�Ȥ(�sӕ"�s�ecj���M�;�H3�yf~K�Au�/?�X9�|U;&����d�� �-��?��k]��ޜ��D�ͩ�u`$����R�PՎ�������T�&��3K#3y��~�m���5<�]�e�M�atب��e����\��Xn*58pY���>�W]�-Nd�Y ���#)�{"��."VV�͛d&~! < 8;��k���#WO��X s�baGn17V��=FW�,@��}�>�! _����B5X�gn[�H���NZc>�ʎ7�װ��Ԃ�q>{����AhXƉ�e��������̄�i�(6)?�vp[�߮�1!��ֈ�����ׯ�`	&�F��o��5�d��b���rdJ�8	���� �T�b�9�#�Ϲ>�C����`FЃ
8����]ne�*������:�XƣC��^X�S���ZQ6�VSd�4ey���j�A��S�r#�G��"p��p�+dY�j���Ƿ�,��J�=���a£�-�+�E��ÃX���
S�)�9o��B�h"�W*���_��F���"!��끠0!�-��Wy�� �I�$qr䙨Fp:�pm��* ��{�w����`��#�ms�L��<eN�c��
�t�~l��Q��� m��9��$C^VQt�����F`�h��(�4gA}O��*Hp'vh+*>�K�D��@^��C�d�+"��3Ϭ����5�O��gm�}�pj�~�K�� ��M?��Y�?Aw`�F�{v���[�_�����nؔ��,�J�Z�!��H�PzϤ��v%\U���R�d�r�Q<���<p\���Hn  ۀ�Z��h�	a�pΣmn��Z��|��(Dg��M�#m�4���@��Y	���z���֕oW�5kD�cbKĳ�[y;f��t��5�(�Z4j��E����Ai��{���,G�k�3@g�'ѳ��ۑ񩉧Ā�!��iM�!<ȩ�䬻�1�j��p�h�<�)�|��R/I6���53O_���
�e-�/��Sr�FK<����
�n�Snh像�����vlV�-P,�(���y��]>���؛�K���%`��;�����=��M�V	���M��Q�����z�2y �4_gI�)  f���G�V?��v���i�d�U v�RI���Isjs0��M����xUYd�ꦩ~��/z�+e��7��F�41{?py�Y�5���vq�����m��-� s��t��B�_>9U�N��nS���-�4��m�?`��*=���A3'�q]�،~�N%3$"��Q��^�C��$+5�i�#o'ƽ1c_n}!�o�z�ɵ�㐳�m`fh�ǁ�:�qL�+,J�@��D�/�' �t)�)(X8�tS��<�a��������`�(�E_=�O�:�Q��]n���G�B�cj;ѐ}S�K )�nmt�Z�2t�%����&c��U(��7��Ig�q�|~�{��o��U�b��E-�[?�^Wę��)E�f@��K8���JB�۾|܏:n�*˩�۸�\'�qʒ���pލ@�9D ��g�i��G�s�$8xxƺ��Q7��ʦ>&�_)�.E���bބŲ��B���c���q�Ք���C���,���5&<��']�I�8ַ��� �oB��S�s^ �.��dw.V(�pۢ"�!����:�{���}�ʺ��y%vt߄�ʗA�g�M_�)E05<�W��zfv����	D�2�����8>�ę���Ό��s�I�ˠ'u�(j�@;��2Y��FK{ߟ�Ԅ�.���J�K�aàG���Ъ����U}M�z�xSb�b���e^�i㴰ҭ^aS~�lqt^��9}Қd���{�@PyV)������(��fU̕��%up�3xj����c�)� �G��b� =�=
�ȯ���~w�>M|�n��nU���w6ٴdm���T�[25�[{��K!.	���4�V�)]�7������/�����6��j
�9�,4D��˂v�M�*��T�\P�;Ԧ����k�G��Z�Һ�dBװl~ӷ��6�]�:$�
�Cs�}�7�<,*��F n�����x2��a���ef��\]���I#g�G{n�Y�6���N��*.��/��]���@}��}��|����2�@fv�ˀ��T=eu�O$���ġ|�f��|�γ����t�)�2���<h��TÑ酞�;���ڌ��ʕ���	@���R��_�n>���>I��f�g��A� d	�}�ɛa�6+�j�=���-�{ӆ�9��!�}�)��{3�sEn;!�6��*K�m��1�J@��jl�⤙L���h��Уp�\������5cu���zQ��*>z}��˥_9�B�g,��[Jv(��¶��j�n(Z��Q�|]�Aԝ��y�e����OnU��V�2z�dV�n�o��jq2d^LީihÊ���'g��@0���3�Z06��R��L�'M!o�(��T�qh$Y#y�2�0V*�ޏ��l{ڤ���/�pd�p�hf�^r-�?��%w����ʆ����P�c;�Mn^�^> �Be&�ک��L`�ܤ�*
��8Xn�;y��lB%�i;���3�5�!9F\�h3�c��Bp%E$ج�=K�$�������I��ֲ;��{�ai�'�H��Iç[DD��H��M���$���Qk�_����~�B�8�_�ͽ=��#@�a�N4yQ�A�<���)k��C2����UwBX�,�7˂�#=�6t�|��H� �9 dC�H�b�G��;��tpp�ojM6��w�'ga��<|�t�6��'MZ��$�/�K����ֹ�>(r�{<�Fl�dI�|�q�W����{k�x��ui�hi��I�Q�&��l+ű⃦cP�����S��r��ʜb����d�3Q�=?�hi�7K�b�Mr�f�e�гN�Bɋ������x�2�/!�t��q����;�x�瘛���Ehڢ�R-�/��Q��q��|I\�%.8(���"CN�Ag}�+����~{�@�k+�y��Դ�N-8���ݭj�5�|���Tn0�H�X��[(NB���j2���?CgK��,�w��n�
ɜ���YdI^<�^��>��ºF��y�o&+=��c�S����9��M�zO� ��Α�@j��tz�mCA�UHac&TAk^Ce��~�H���zCW�윹g�β.��,#�mɳ�Xm2��y���F�/��t ?6O����%�ͭ�fR���ʨ��Q}���G��C�ֻ�9�cM���s����hexjZPmHM��r�ˠ��S��� ԍ>�Gx��eS�=���U%��w�8�jC@����;���1�����#�P�H�Tc���!�:=ͅGZ�P?�:pq�ϟ��Ԩ/4�hĄ!�B��dm�/99)Z̡OJ�P��n�}������4���;:�ػu�p��:��N�58�,�����φ��vq�u$ٯh���>� ݄[�� �ͮbi �.Tf!Dd�Z�z���D�5�O�`��.�a���@������J�����[X 0#D7�`	��k ��^e��@ZM����(�ͅ�E5�{��3"V�4�~�d�;��+t�O�g?#��g�.�a,�!G2�7��Јm.��DqH
F�H5u��$�A6����]�-�K�Ѵ��d5�F�׬K��{;Sz]A�q�ϲ�\GR2����V`Ǥ�EiT��I������΅�����ꦓ�b\�����?�6��J�,� `�@�(z� ��O�_�s7&���
ލT�7)5j�����9�*��<�Bg���P��W$[���f��%Y5��2������ׅ1aXuW���aY���U��kBr���̚���O����+�O�yq����A���{���x�n�t4����A��̈�Dү�	Po�Vب�]��pU���6H��))AT� �I?��̬&�;U/"/�:�.������YAټ�����߹�sA�*�9�kx��M�#o��OdZ*
����<�;g28�"���y��R><�ա-2�Զ[]��5ir��/� ���A���S��n[�C�w�^q�|���(�u��a�U�g�J��
䬧���"�'�f�-�6����pk|��2gkl�Z�8<�H���ݻK���ʅ�#��2𐠛7FBM���=�t��9�*п&0��$�d��85!E��D�-�!��� �Wl�3�	�}?�B�������*o��w�]�O7Gmja�V�j<uL�f����<�jv�J,���Bm�&�?^���v_��մ@}��=�f⅙/꙽T�QQ ����	L�L���,��0^��6˒�uRl�/�o1;{,�6��!r�� �@v�)���>�z�`�H~�� ��[m؅��r�xX�j����t r�P�}��k
\0�0�m�����+�Gm�>:�cY�c<�2��:�i�����Ng�VmU�R��E&�����N��NL���s���Ie���;�5�u�CՏ��g�ፁ�Za�)O#g%˚�n�h�����A�6@���U�Ck�:j	,'���V|k��V�;X��V�KY��,��gZR�.	�^�����'f-�Ry:1<=��"�|g�B\�l6&��(���1jVI��aBxj���kgx�dy߉ϮT���<"�m��>��}��Y;��X[�����r�(��)lW�*Q�W�QRi0�,#��^��!�=��t�ySIă��3�#+Q��M~�S&�EC�j������Jݼ����,��*LY�G2�7Q�a����@�A�z�k-�����O�ܰ5�ñַv$�}�3��c���V`�;���ED�`-�sBP�����cA�c��N���D�*w.]��x�DQ�͉��c��E��!�M\�����D���&[u�H��WTTd^�0]�1)��
Fm"->yU������S��o4��)�s�J���(�]J��fU�^���s �u�چoNy��1�(h���,�ێ�ݖ�H�� kuj��m�Y(D��e]�r�P����ܥ��n��*�r���/IZ/(§[��Iy���r�����Z�(H9�	^�LY�H��]��>�H�x���#�M��S�v�q�1:w�lZ3"��SV0XI��tɾ�yk�C��[3�
q|��a�{Xa���A�� X���la�>��M� �+o�u�*��^�ecCHM̭��������LN���,*0�`h}��h�NC�5���q���ts>| Y��pS�8��}�\sʆ�k9�|�t�%B�NhI�MT�KیאR'ou��{�k���
Q$�b�M���2Vq��������838�D��v/�`�p����L���DI�z�nb!�z�焍_.-R�BN��_�X���y��߬_}�In0�.ʫ� bUpŢ�m+�R!�.�g�����"��M�)v��<i;�J�6*K^�������K�[e7pK���X�]�L��n�E�0�v�ljt�M���j����2T#���m��?��**�[W֚��&�"彦6쒝���\������p5�OOp*`s[�y�%��G�^i�u7�l#6�i�Di֝ �bf~���7Q@�Q��W�yW�>#4/�[�N���/H	�)���)��]�۔��;M���js�s�*{.F<�L'��ߐʩU!|��+��B:���������Y�:P��t�)T2)"Cٴ����� \H\��8V��;�����ճf���n��?PU��R=k����Y�J��;�G����o#�4�Xγ8r[q�&���֝��d7&b�
��y�&��T��_���1�4i,��Z�e�%�����l���,�@���g��8�O��Խ����j�n��~R;,�`�f�.Iԗg�	n5�;�>�=0����AP��h��t��4�=!Au�:�ۈ��p�t�(wt�Ѵ�r$؟�:����w� ��A���Ip#�h���:i�A�#�>(���lng��?�S�0�
��eN�ȶ8$���|�����a��Po'b�©�&�~1��k�QR�j?@�J���A��_�S�a�(N��O�N>3iv�Fŭ��������D5 ���M��^�"���`{F
N�%+nC�ʤ� ��*���Ԛ�
ó��d���Ҹ�$�\iz�.c���GghPl� ����)5�,E��q�İI`l�=C�E��;�IrM:�w��wz��Y�M�ʵ��W�7��NQ�ti�Z��q�o@�s�bý�;F޼�P	 �W���ϲ�ҳ���:Ț��o$�m8�H�8�߈NwU�EK��k8 �(�aS)�`%�b�\��A����EasOb����E�E� �(
Qæth�:�����j]��R��I<�O?0��Q�a=�`���$���*�����u��Y��ƿ�� P�w�S_U��^ƼrH� $3�.)�
I�5|�IGq�bR�J4T��s��z�G�7sq=�.��s\n�\j�����1���S6���&��!8;�]c<K��>{/�C$��o�Y�D���7`Kt=�b"�K_ȁ�f�m��lD��o�7&1r�!u������|�ҿ���3_�PҒ��a�}��)�ⅼFL.1A=�O#��!�n{T�Ϧ�w&�W�e�"���T|�פo�/�:|E�oOv�e6+��7��l�r5̳\ж�޸���"l��n���V%����99�fz"GЅ��`�mv(���7:e	�0�ZY������֚�ئ��q���3�h�< L�q�#Fz�<��F��4�?��7�WIN&,"�h�?!����#�KV���l��.�auG��}�?L9��8p�1�:����Z��������&��w�F�0�g�N�)�W�;�v�ݐ99Et�]J�u5V�"�n�=�IJG��Ü2�'	��t.'"��"�cH�Aʋq"V `�D�ߨ}�*��[UB76�,`6��4Q���9��g���)ܒ#۰�ۥ��G�q�M5���_Y��7g�BQ1�P�a�T.c�������*I_���fr0.�ބ"��#`m����$"���UR+��Kv�(���9����~�Pri�P���5^�l`.���A�(���1�����V�J��+k����yp�- �������dEa����8���ٵ�S8j�(�)��F��Q�+b�����0_$R�T܁��Q.��Kll�<h��|��6�Ui�H��߯-�=M��.�1���3�7�KuԺiѝ�_�D�;�-J�l/�즛��7.�6��j?Q��&���[$yZ1��Ck�b6h�`�܋�g�|:����
s���n�Q3�Ḛ��ЏAN
��b�@��R~��v exd?�*� �3�CJJ ���Ǽ݊T�~�Lϲt�=s�^�A@���´�������X�R�\�~5x��׹{�I����<�NbM�N#�����R�Q+�<Z��
5�s|[�Kު(0�E����&��Mљvn}�ٱ!�Q����_��ٕ�ͪ��̧_����������ȒT�G���O�g}�s63W���[oP
'՞}oX�����1E޴������{n�@� �P��y�U���(8�]��
/��6s���@�Gk�&��w6��J���:uNs&������zjt�iM����8.������vХīe	dP����"�=#��o,X�ٜ�i�o����͐��EQ�����'���e�#B�?|�]R5V���x7��	������]�W^W�On�`� mm��n?��K���w�U�Ղ.S�i�|+����I�ki���qd^ނ�E�8/�L��&k'>��8��E����7֖��\es��祓2�^	*' \�-6�~���t�(��ٹY6����f�70x\%�a���w�C(Q�A��cҗ˥m�Y1j��Ox!%0��0N������[�J��o#��������U��#j(�N���J�Zj��Od���M��M�]�����ƙ���g#���E��kr����$���$�{H�.��Rn4j2���s_ P�g���zw�]����Lu�=�/e�4	��Ș#h�0��?�^�LV�w>�>/h�) ˢ�I?�S�Z��]j�
H_r�^�p|�:�E=�W\ Ӹ���ꀽE^�r��?l� ��үе�c��G[űn���?�k]�\�Xz��4#i9Bȡ�{�t��M�u�����0���~��SZ���}�K���ع�È)#��s�k�|����M~�O$�
骕C����0U�c����)�� G��J5�H�<t�UN�V���IQ{V(��^��~+��Ŀ����FjRp��f��w�km�+�(��)���S5�F��o�S[2<�nA9j�N�S2@�2���P�S�Jyѷ2j?�Rp΀wa��ET���84��.� U����{��Q/W�o�Xĸ�/:hp���g ���rc��g�Xc؜;�w�M�0�-�2EBZ��
	h��`M�m���=�a�_cɑ.~2�X� �oi�U�c7�4,=�3���K��>z���9'=;jb��,~�����Uy?C��z��[�<S��f
P'U�$��P��t
�.���'��p�{u�YB�h3"q��Kq��Zeϰ}���,e���Ĩ��Tn��E�?�!a�[F`}6�TSx����6��HB��؞�2)O�;-��)5���}����Po5k�(�]�@?�N*�rrn��_n�����l12�_�Ӏ�A@
�%p�?��Hi|&B\����L<h���L�-΋*b_�ؚK��ØՋ�ɋ�
�6֜+��^�����M&�>.�����B�}�ps�l1������&��Ix\��T�X}��(� �ڞJ:�{g��~Ew\#�Oq�R��+�{�ﯘz�m�%垣�s�Me#�N�y�A��CMnPt��*f�DX���S�v@�s,C���4�U��ck���J�eZ����(8u$�ڀ�Rn�gX�L�Q-ߛ�'�w�B(�� ���[���حj4���33��d|�L����|Yc5�kh������	���Z 
"�%
���N�L�l�U\��8-T�I�a�h<p��y��b�W$��KK�N�+\Am�1�;�ӫ3�&0���Qq�����8�`"y�t�����?^�"��OtI\>�������R��e�:�A�t$����:������k�Ws����V�`u�R�Z�h�!����
�����&��r0tu�������� ��<��ʖ��#��;�UIM��}�&���0],�<Z~>վ��*e�f��A��f��s��zI]�Z�Qh�t��Ů���!:�o�4r���Ih��xº�"P��O�2���[��b�2�`unK\Osk��KI���A�TI���QP��>I��<��NFP�
����gClg�ƹ�_�Bnu�`r�j�S
z}9�!������JK�&�M1��	+�et��qYOv�X��?N�� f���$O�ЌLʬ�Ӆ��w�. ����洫k�r@2���M�$4F�y�[J��e��Pa��oA_hq�P)�*���'�Z���cfY�q0�xtМ'�(���KT� Qmo��S��o��"ԟXbM�L?�G�[X��gθ�%��������ԣ����$%X�����T�?�x?���w;�q#�wl�t3�C��\�	K�s�O�;�4���+����l��w�h.���_$sD;@����	�\kaYb#��C�����mb�V(�ħ�B<}����v]k!�=���`K�M�|*/�E��>0�y� ��=	�'��{b��#'�=��.23Lp��fs$�n/_���Э�A��sD����$m@룇��x�X݆��q��g�,��}�ZZ�R���n��3^��f���	ƪu6���{���m�<���O.�M�K ����ں	�Ҭ�<��eb���%R��i)\����2pDa�P�zC;eu�/�Z#gN�5�*�!���E��V5�e� .��ף��7/�)c��t�pC��z� Ѽ�x��Z� �^^�!�o��&4�������3����9�C��ᮜ*~�<E�^[B/�&�&����y�b�RsP��#*��K�p�t��|\Swv�M��ܹBxg&��B�Z��H��5>i

7ǎ���E��`�H:���N%uI�B#��v��s�f��:U������.�S�izCX"��v$G�W*l�"�m1�4���C�;��$������)�;׈c�Ӿ�q�A��)�*&R׸�T����z���'�r��-�:A��4EVH�cQ����/(@ԣ
-	ǥ�9#�+b��^l	rJw�&�MLvʅ��W*74qY4�hp{�N,T�71�m�,$���@�w����NN첶�i�l�N�����p-a���VY�	�Uc_A�b��v���p٘�6P���N��4�D��8�!������"r�b��S�	�ۚ��c��9|�N�.��A�WFyF�(FhS���P�"��� ����Q�l���,�9Q0�4Rn����cV�)�)#�J�7�۷����	=yЇ
�i!�*�{�@z�ŚI�0К>���3�mWjX��M+��;|���g���-�{���-ށ�L�O��"m��[.���E���<����ת>���**-��)�����b	���u��n�a}	����BEBB��/�nB�9U~� ��	B�L�9LaJMO�CB�6�s��r=��K7��5k�iU͹�,2L#g�ɕ�����=����M�i|���u�rd�@EI�S�~�A��dL�ߧ@
�j%�5���;R���V3��[���K�ڣu��`��d=W�&�gU���r���u�����s�TY��݅2��G�<��`��DTH@3��'�����T�������i��Q�+Qk����`r��wt�|Ϳ��.B�<���gՅ�!cJ��eޝv���HSe�J6�E�$5l|3�k��ӓ�nk��}�^���V�r핶�h�ӏ����vV{ҍ�z����+�.IH�����]��R��m3L�^9�
9�
HID#�{뇢�C�d�LX^���h'!��T�E���u,/n̓I���Lor�{nQ��Y_|�g��'u�O�����$�����0�`Ђ�_�٩|c	�46H�	{�`�aDI�ז���"F$)HC��|��ci1�.}��B�Ȳ6�T���T�e���(ǡ������\���O=�5�[{h�N������>��[s�e!O��S��a	��f����:��y�'�v��_��G�:t�"���C���0��a�=��r�2?4Fmj`���#�.P-�9M���vM�G���ɭ��3�X}ڰyh �K}�����:k���8�`i����!T�Tߞ���0��1�����m0�7��Nݓɤ�;m�)<x�V��ZY�����D8�P~�[�50�� ��it95I�%�
�`����t��^��1
2GY�w��# A�V�K#��W����r�~r����.���<J��P��4�4�ݬ���N�}f�Nmc��J�>ў$�d}M���I*����IPl����@������~RA��Q$�{�V�@�-R�:P��='��P�!�G�Cjm{�A�F�}S��~	��.�w��[n_�#s5�A�$t��sjv�[Pץ��I�1��_4����;����¥4�>������˻^A2����t֮���D�x���۩Q`+�1�Gր�9�徭�g��f6Nf$���I-5�qD����W��������c�6�ޱ�7��G,�s��,J��n�7s�@��\�����X�Y.`���U ��o��Ŗ!��mv���$-J~�S�p7su���=�|���I:7ʞ�`�=�d��u��u��/ir� o0!?yV���0���wl���6�K)�#�wp�yP�%肰G����I"�͊91DTqݕ�҅ �ra���w���u��p<(�A[r�"����3��'��} �HFX1H�%�4���>�*�OvGd��[9@x{lZX0ժ� �a���w�����I��ϑN��/稜����*� 1yV��t�,���썹W�W����a����Q��i��H3�lt�)\E�x<c����߬|ҝ�`D��߬�b�
�m�	Twa�6��>�[��f_�]ė��颓��h�����Q~�#.�AܠL���7Hb�+���mp��������Q�}ڈ�����W��������_�]S�����w���)fE	~[�8�&uz*e�4�u��>Ο��_�)3�����BO{��plGH�3g��Kw˻AK)!�� 5�Z�qz;�5���F���] ��;R
���н��#��4@�?�>�-����s9�h�{5�QK�t-�H��X�?��K䡱�tl������K@go�zn�Β�K_#��z#�Р���<T�/�2܌tb�;�Q�B�|U��[,i��E�l0*����V�hlEt�'�1l�x��DF\�٦��Js.��Ț+���'9a(0�c")Rw��
��Ɗi;��/W�=��S������&�w�������D�|Y��n�ќ���(�J��*��$���e��O9l�vT! ���rN����C$�$>�D|V@�K�`��N���'K<����
KIӿ5>��F��#ǽ;�b��[%�p�d��H�NjfF�_!nN�^s�6�+Cp��~����#���Q[%L���m@�1���W<��9(5�GU�<Q����'\l_̝�亼2#���L��%�^e]L$�=��NDG��x�y��(.o4{�F���
��� ?0����9��U�S�r��N��-��-t����c���H(v�#���k����>��C	"9��-����c9N8�*�������4���.:��Pڋ`i����휾3�P�4(t%8dg��a��9��`B���_�w�7ӆ1d���m�1-W&J)�d+L����Jn�.�(��1��#n,5��-��r��	$���pe{�+4�T� {"�T����L3up��(Q���p+�E��6�#?�O�	[>�m�~����ܯh������8%�t��F�m/>��E^lr�uR�}��em�븽��ɭP
�5�{�@��l���S{�2?��ίl��9���;VYN�ȁ�$kIc����li��Ye^�i�e0Y�M=3v�N�9>�G+
.
KZ�V�_�Pil��|����es_�ğ�<;�J��ο(��З������nW�@�#- s.HJ?��{�n�&X{I�G�����O��CG����)�s�G��S��,N�&&{dz���'����%����_Qm����J���XC#d�;����ަl�Ę�U`��&r2S��0�2Q��3����l��O<ś�Ɂ�|�����T%����8���q��� �r
�pK#�Xh��\z'����.���?STe5��@������
��֍<���!Ǟ۹�M�+ �5�4�-!��>Xk5�ع�.dX��	�*�4� ƅ|�'hU�yg�8��;<Ȕ�e��^|;�e(vA��J�C�Oh�����1� ټ[���;��Ũ1�L8��ȳ��6��A���&lH���:e\�Z5ˋ�{�0#tAsR�vɅ��p�;^��~���1�<	mb
恜e�D�ѐ4[���$Gى����`Gm�]�@�S�XnT�YP�H��JW��%��\V�F���pr1�����A`������b6Jt,F\@��?]�1p�,�c/?�S뉱ā����ւ�ZYAo#�<d�Q���
Z��ˋ�]u\���Үb�#%�&Iܝ-�P^�5<!�+��'G���x�h*�z{ŚHl���x;����U˩��������AW.q#YL�sf��qK��F���8�nU��t.��f�7O6\�FP-��b���{$��9 3���2����ت�RS����we�L~�����}75(��V�� �E��;�U#J>�P%}j�BSM��p�E�@�(����F���Ud�8��M�N���Pf�Dg|�~7�T�V$�g�Lxj�l9����ׁQ?�Q��`$��q�g�b�+u$a���wT��zC�_j1m��#�J��G��W�\�en�����ЪsIM���7�����sn�D�k25����t̋�ux�AL�|�^������W/Ĥ����%�9��DQ�����_��Y���}��gB}��;D��M�H`[��b���t�T��_A~/ �3,QQ��+���w�pb��.��߫u!-�b����^Kq���J hC.C��\�mUt�w�������_������c�hO�d�KJ�>�q+Z堷�.mO�81 ���y!�!�ɠ���J%�J^�uy4�~?j8���gH�I�����.|CX	�!��+��Ca�m�e1,TI��\u��z��8����en��I��ᓏ�T�g���[�� ��\%��rVO����� �f��i~����~1�Qa��I��O_�o��B|��3���󏁀���V�&���F[I�
ȭ
�J!g�gߒ�P��[NFjU��.�������Y��c����~�q�`��0�~F����U��,!�޵,YDo�8hQ-8�& p\�X.}��o��2]}F�s ��Z}���m�/Ui�<k�.�/c[���S�r	�rV&�蚝�(^�QWw������팙+r�_���9"�ڒ�t0OL" ��:y}0�Tt���j�h�������@/OTF�L�iSrR�
Ƌj벶M�ʬx�L�o{o?/�������C]W�������'j�1R���AXe�\v��l^��mHw�s��y���$�ԁ���oRp��;�D��/oe�v����%�W���a�j?8F����Ǯ�m]gUɜQ��B2q�z�;U�ڛ�]����ᘫ6H�������l���	���%�)��n�_L������H��r~�/�J�>�`*4��b9�	x:�Ev�ٗs�}M��>r&a�#i��5p���'#��hl���-;J��W4�~�oN�H�5��qzvY�.,�MW��:�MGD��8�I,����62:���w���!�|��q��{�d}U3�b>�&VIk��`
��6.�ÞΩ*��b"N��@�IX,�� W��vu[Q�����@8Qw�(�Ĵ�b�
��@2�V_�7BG�;�2��`x����P�~Z`��&��)�uI��ǧ�G�
74��6&R�N�6e�B���P�H�Y�wǶ��ɻ���@��rܚ�;l�l޿�]L ��t����_�>�hoE�b�ʯ�	����ܝ����FQ�~��$���t�^��D�۶TV��g�TN�"�gm٨Rﾏt4�hM����+�Z ��
2��"1�羦]��vW�J(��-� $�>�\ɚ��Ls�z,4z�Ă��jB�_y���ID!��!8� !���=V��RTSD��֐�Y�H���H��R��a��$��#��d.�ݼZ(g4��3��6�%U鼼Y����E�>�?K���!�JmW���V�ǩ �ȁ:\�"����������5�k�'�8T;ֈ]đ
"R��S���<��0��-s�	@ЂDԩ������H_����x#!�����c|�MK��D>��X�-rrx���!nPr̘X����F��Y�'�� ��Q���-/9��a�wE2Ƴ1��x�V5scP�*j��d)����0�(!���~�S�V E����,Tg5Z�.�@yx%�p�7Г�2Zr�q�#`X	Y#�0�lw��!���M��/zՃT0�^�ޱ�Vn9|���hxԤ5�J�c}�q(+�&Е	�	(DAd����-�F$m@0n"��=���`���u4��Kq�l��O�6�hT�	����Ԓ��\Ye���=��5r�,7���2Ұ'!�z?X�W弚�E=���k�"ݿz�d�=�/�z�˰�yg�(P��Y-�>S�/n;���d�{�6p�2��z<��}�㎫i��a�<9t^��s��%ru�~�	p�JW\\EóLT�?s\0;v�W� ��v�^�T�f�w4b�Đ(
m~d��H��Qd[d���p��b�5"�.�d�Q?Ѱ���Q�Б3+��6���rE�,�)3����|�r��4���ڦ��@����Li3
��T0�[߭'ΫA9����V����W���Q\>1��u�i�!c���x�4F������(*���K̠eYΊs4��'��'���9���2k�M}�G�i�K�Q��2b�;L�8i/�����٨(�L��t�g��Y��1���<gD����Cb?=+i�3"�NR>�TǔtKx嵝�>(��hr0{܆m�n�3e���Ni����Es	����ËG�3�#18z,~����̢B}�+
:��g2�:ʻR���b��P�O�����o�p;Aa�!�5</�ͮ<����O��g�jV=�B�*u!@���2|z�R6�=�v&D����h�i�kt3���j k@�Ɂ�=�>k��>�1�z|Bb���t���y�m�0$���)���f��o�
��P�O�K�U�ؑw�+9�J�O�~Z��Lt-h�I�����'Æ3Ѥ�q�K��/��wx�- �;K��z;GѼ}�h��R�PP�)�Ź\Z芳K��>>���V��Y�t�~�M�O����THFz���+��(�H�HQM��i�_;Ἔ��~k>~��z�^m�0@���J�{�aֺ���
��G����,+[dnڄI5+��l��:�e�����.i���{�%�M�=��A�?�Ȉ#��y�і���H�m�_Л>���N��V=���m5�a�!m����-�^� qk+)���������Z+�@���2���2M�8�*Y�D�(?5*�C�������|�\�K&�"�a}�U1�Z�'���7�����f�eM]-Ǘ�3G�C�a�~�?J���b�]ϊ����@���ӑ1���ٟkaQ�M�diln-f�Ë^d�|� �t\g苨/�����'/��(ΐ�G�쌷�|�q!k9��x���ALNp�W�*IG`�2\'��%�����Е��$��������K���ض�l,���_H������ʩ]��m9�P��t(� x����s�g�g�挤����^,����=dNfp͕�M2�P�p�]���:�T��LR~�
u���mDa����4,���� m�T�|*&�As%V�T[-���3�@�*�EG����Js�x�h.6:���OT2f�WuO<Q���aH���d�Jk�E�\f��;��R�w��O��h�a��?(&Ŕ[qz&��_���྽���5�W��,�]�C�n����g	@��o�(7�]����ގ)x�)�_���N�n?�>唀2h��G��IB���Zq[��-"+*���;�AE����h��EII~
�o/�@|]�� �߱S|�濚����H�;��(l��	�2׿��Ы���U��f��4�L<d��Bj�԰���o�N�b=g Z+��\J����^�8��X�w�ؿ(]��y	�m}r�4�2j����U����N?�n�ka�c	��h�.(��>�/b ]�v*�R6���l����Yv*�Ig@]��-��p�A8C�a�La~I����Y^"�,Ҿhņ&*NeZ
�E���{�J�B�.�S�Iu�x���u{ h�),�ơ�7�8ߘ+�F��	dd�����	_�햹dÜ�r9Z�5�E�Lu���|��c�_���9�����!��RZL�
��3&�e�+@���:�b��pm���g+�h�y�՛,�/�Iź�|.�k3��6�>�6U��1E<��P�8���i��
�&@.��=}ꄡ��V�VtX�woJ�!TYqhiz��<��zY�G�f`u,��1���*���c�Ok.������E�;$��i�o�p0�V����ŞC0�kc%���1��<���A�~�`��D���φT��k- �&_f-ӷG��_#C�Q���6\��_h�������`��T��v-\n6磡P��6�"�7�S�.@���2e�z�ܚA���[�B,)V��\�2E� ��2�b)��峸:'�:/��|��B׳��ԓ���\MYZ��D>;s s�������Oɭ�|\f��_0�Ѫ*�����K9Y�ڮ�����/�.�������t��>�ŉ+/Jɞa�x���~�Iq�v��пg>g�w������g|��39i�/�D���E��므z��L�w������ hI,�n��r�H� �f"
%j�9phԨ�}��h��frzj/��)	��v��7��Fr�z��O�Wlvm�߈�)#����C���Z��V������p�Tt�U��"��V�K䐛�	Y&��aT���½G$j� �⪁[+o�@	feRq����ʻ@�g	�n!f�Pj�}k&��耬�!���_�je��4#���57Igl�ͩ�ғQQԤJ�1�~V�?�i	��(�i�W��.��(�����6Q���[�8����^&V��ܯ�Qj61B��dXU>=��g_��2���r /bIn�$�Ҟ{�Ɲ�5�R��	�Dҿc���r��3�z65C�]jaP�B5�4�f�f��D5��60s{�N?hK���4�_*��l�m&��dWJ�y<H��U~��{��op}=��I��~r�����_Mb �)�W?>��޴q �]U����Ҫ�)�W_*`ߐϠ������R+�yEB��(v]���hP�ߺ\��)S�K�&Ð�l?>���a�S'k�%J�(M��Z�ɡ���i� H�aܡ^-W�q?�� �vx��쎶��Ư���0�Y��?�dQ"�(��oFIz���H`Y�Lq^~�vu3\���tO5c�}F��w#�\��i,���,�3~��蔀h��ma�*oy�V��zb�cdW�����	½�A���jWF8�L�V-(U-D羽�$H��r����铝���Z�{	J�3""���׌z�6���)컩k���R�r�iF�P���ϱ7�J
��f²���a5���e3-l��4��+��'����B~��PK_�����X0�� q�勩(����pβ�����tΘVw�F^�ts�"������%H
j��B���|H\�&�0�O)xɜˍ��0��Yi�N̙�A<2;�Ռ�|�j���<�~��zL�?��O�)�*8��؉\&MOś_t;{7�A o�]<Z��^|����g���0�X)�6~)�;i��5�?�$�į/B��H��#��fe��r�Bv�����"��a8���k�Q���b�>*����~ݩ�'G��	 κy��'�JVu��s�~qE�l�:9@���o�����_ˀ��G���ib������G?����{�,��99��'Hx��ɩ �Í#?1Cb+B���寉P�4�L�����#x^������l��X�"\)��b�TYJ���;�Ú�O��]M���-|�_o)=B���ߌ"�b�M?�#�;�LC����o��N�Zf+y�A/Y�MK�\��Π�+;H�~���1�Zv�W(���P�C���;��5W�/�S~!}&�m�EV�B ����빇���-=���jVQY35�X?����B���ª59�v6�?ؙ#�1БQ�D5��Q%+-���D䕏8�����<�aٹF��??��fN�'�Gc'��Ԫ�7���� �X�(<�!�G�o X��9����{1�	�w� ���(��)�y3��ĒLј�b�������E�E	%�w��{������� ?v#�q�P/�&(��ܣr�s=/�i���P��H�d81�X�b�gx�6tN\a�������(.�Y~��Q��l���=��:i��wf��������@x�H-�a�}�u�?���R$������b��Γ|����-�s�A]��i2�1��F�:��Y�\���I�ѝ�f��<9x�$�zPp�(�\����	��o��͖�f��kLP�R�������E!�.��K�Ir��Wj��K�>D�d�9P����^c�gR'H$!�Tm}����,��YS�vK�׸ g���]ەxM���'�FJ>�')O��w����G��h�@'���Hqf���Y7������s�b���e=i�;����'�{1�p:�I>���p@ v�����8=`��.�����)�E��>�w[���}���Y��G�">c��UӁ�h}�2v�F_jS4��Z���)/�u���`i��ל����W�?���]�<?��K����l�h�9/�F��J�־��D�R(������(*a�>~����Jv�U1�����f��ѡ�2>���iG]@E�O@�V�����ݤ�"��"���myH Ŕk�4�P��8{���#n_!�<~�l�t�x$���6�����K]�wǩ�!�^�0���1�Ĕα�zXdpÄ���������S舠�tK\Ģ�*�j7\ٓ�g0 "p�*��p���B �J�9�]֢F��ԋ#�x�&2ԛ�H���W�+�H���Ɋ��i,�C� $���2�8����"�?m���J#���|\60�7V/~�Ѻ�D^a�C����Nh��9�M�c��O��y0�1��C��!�L�פ�4�`��ԗ�в��\9qD)#K�>�@j��8R��-��^�J�0`����ZOȯ��4�uU���1�~Y�?x�{��\#�A��0�)t��|넭���9��*E7죑Ml��w|A8$�W��H�cC��ܖ:�eE�俞"��2f����uM�^nSӄ�=��;�����W����&l�'M���_0��J�����"H��E�ҳ3�^SmAi�Ov�1��+�"�� {��>Њ?O�������c�����%~����%(�$�����WЋL�Mi]��~������=�b���,|*��<��~J^P�4Qi'�OE���O�h�����_�������<�x��Ԣ�-�l܉���Ǐ��T���f?@����Ёƫ���U� �m�.��1�OޛP���4m{݉�Rl�,����v�4��!��/%�$;��bdi�y{{>�wB�;�W�[�EЁ]P�n�a):�j؍&D��(8GZ`a����%�>w�	�k��怭�4�BQ���M4=����M�N/L���R]p/ -T�قϺhd�����fi(��s�k��J��)h��r�&�A<B�ik�RC0���N� ������蠆����a�J�M4ը�?�z����`ΘVg�vflABpb�k�G�xhA�E1ߊ�����"���IU�b�X��Ő�kO��ȳS�j�ng�L;C�R޻�Q8��6��y�8���AѪ��չr����-���4d�m��U 8�E,�����N;�(���yڧ�Z�
3��Is�п��('�{�aB�Mk����J%��Cǣ��!�3Ve�حz!�]48,����T���������gjޫ@E���aQ� ��`1'��U9.!�#t�A��4P}�ͤd�Il�+w���ɖ��K�n5�� �v 9=�I�_����)�5d���/'Ǌ����'��~W��9[sw$uY�J��NcxqDK���S�T3��X�$=J��饬fIM�G�g�V�W�Ԛ��4Iv=��ƺ�MU�@M��S^d9�{��ܐ�TZ��]&�ٶ-�o�G���e\�t�� B*�4�~��+=ͩ�����la/���'�dM��*~ޭֶ������Y�N����@��6�΃%\-���R�sfЎf�z��������2 ֘��<����-�*���I.��C��t{�4ò�o�K�����ذ�	�����ʫ`4��"�� Gʩ+Jd`��옏����|�[�H�`.2O=i��Z��g�b�_��:�Qj�B��p|~1g�����h�_�`�+e�=��{߰��l��KZ���$6乱ʥ���6��4��<�T^Ƞ~/�&cPi�&`cn���-8dd�������wʹ�G}�[L����L�Z6T:��g����V��>�b��,�S��/ /D�ZI(M�fz����=*�!P��	(N
�G�/»!e~�!~���)gy�D!�j�Cf #�o_[|g�9|N�95E&�_T=I�]��D���0��B�(�҆� _c��yc'�T����~��1m,6Ό�9HD����O�ϣY��b�P+�(��E��������i�Sq�(��Hq�K�[G}��X�U�=�*����wm�!ĩ�.����0��1�b	A�K�׬E�4�o��S�{٤ He�DN߾�+o�o3PC�=	�+�G��h%��{+�-	;���~�R-�S�*||]<�ҏ1;U��(�H%�,M�.r����8ڧӰ��:~����vM���"ۨ=��S���:Qt^�9a�\�Ȏ���l;XҼ�]H��2����ʔPv&�{�cn|+/��YR�\�U��u�A�҆l�ļ�g-a�-+W��Օ���/2��r�p�o����	&.�q�ոl�F�Ơ�x��gb�s�Dk"�$\�v{G��U�k{�6=t���7q�L�yV�aDN�oT$;�Н���H@X�i �_Rr�䩎�Ր[�l���T����9������� �T�WN��GT���K���ma^��/l��o~�6�){}����ۀ4��O'@ �)g���}��H�B�E�ۭ"e�g9�I��6y���@��xk%kM1���ڨ�5 0-�?}�X���kag�
	I`���~]�A%��%��]��A�u�L���;C_͉�)�c%�gaM��o2m�wE�3H�)c�.�����[<e[��L�p����HCXݡ��Գ��k���M��ؙS�ܚ�ۗ���pL�L�36��������D�W�O�R'���#3jA�y�����f��a-������a�2Z/{�*4���1r��Q H3r*���N�ڬYh�xL�728^����8������Z�D@Uw��#?=F+�#�g�~��N��ǟ��C�kf�j�:{}]-F�?k�=P���81�AY�����Ğ{�^�����ɾ�e�9jf6��mP��0��8�䩿�|�j6��ѳu n��z��^��:q���w<U���{�TԖ�Z�j����l0�����y;�s�A(�ϴ�1y��@�������V�$خ��5�N�<J��6p*�~1��%U��5�;�0^B�	���x�u��G�������v�R�$�i�V)��hº)���w��5��u��w�����(�*��J�)��	�@X�l)�)�1��:�-�较���������!�*����f����"�6�ڧ#Zy�*lE��yYO�t�u�p,?@��8�1˰$�O�}8v�|�tu�1�h�l!zbZ��}V�	F���*�+�c�k�h�{�J�H�t�`�I��Y��!I}��X�Fvo_2R�.�����[8�BN�ڃkg���p�����l׼���P�hՍ�,N4Ͱ��!Y�)�p����ΐL����4��t�>>��(�����lW9�Ky��᪉����2��+w\���3oV�Q
��ƺ�\�Vi��owHl��<=��w�|�P�#��3O�(#�0�QI�gk��")@=���B{ĕ:�� �0��X`p�q�xk�3�a���ɐ+����m��7{�>D�W���K�a	Jt^�����!��b	"tr����#�~-]}���`G]^����G��l�>1�&��D`d�	�x�PLG�ʰN�&��5a���&]h��m�*�+_=sy+�[�Z�XK'���%k��@#w�!� ��cN2a�x�1w>'_��BO�ߢ��d.�F���HAc��RO������|�ӥo?ZM����g��$��#CK�����8�S�����}a���섍9pH��͍:��P��2�+��P(��
����rZ�q��o����jor��5�:�����ِ��}`�٫�� ��4D�_p(R���K�������7���C[k���%������w�YE�}(#q�����/�l�9o2ɼaJ�R���%�{�/�hn�놁p�s��/Xz�91��Hp�Ikԭ=�ԙ<��3��9�����;9�E}�X۹.��:R�Ŋ6�w{d����ǰ|�R�\jG���ݴ\a��߫��J�n�s����7�f 	���7���ڣN�g7
p4w��ꚢ�=�� ;�To���lUN��lN��i�d�5Q8�$�#*��Gߒo����л��`j����M�����}2M�95�x�U~��x?� *�˕��� N�Vk�Pp�۞vA���6�+qHu�5�]��;Z-�3��r�TC��-דu�(�X�'�T����z0U-����x;�����|=8��B7�����XE�^y� �%�	���c��'��S"��#|l��@$��6�y�<0I�z�� T}V�̙�$݉!%���L��d���ڻu�A�=3�|�����h���0z����oR��눂����|��҂��|��q�ؖ���B���ۊ~0(ѻ1�!_Q�$�MF��1A�q�:�U+��sW�˧����OR%�[J|��u�D�PI�w����'cղ+��#J��\���-�$�GeB��͞O��V�%k}����C�K�Ψg�v�~�P��鋂�2i�EsM
��c���3k��S�0�7f�'(�c���gƪ�mF�_Y��Ԕ��{�p��z�9�l�j[��7��wr�P9���W����ϼ7�M9���?������F��Q~Ι)^�5�������I�W!u��<��W]�|�n�XǏ��8�E~p��}?vs�,J��o
e��'��x��3���<�ݲN��i��'�<��R���-����4ɻ�e�/�y�r���R��F�)7V�����Xj�Ȼ�&xo]K[f>��il������Î3�n�l�!1Xa�B'ϰn�g�$�?ľ��N�O�ݯ~r�ݡA:��J��H��<�J.0V"�_�a�+?�fj�;(��.�~,��d�^���~,�=�;�D�@HU :�?ՏD�4�L�=��i#�	Г.�+���ۙ!+���@g2m���!g��k��OJ��fk�C�av`2P�9>�@�)U���S����o-ɔ׾	��fG�����9!ǝ�U�#;��"#%��ϰX����⧮�c��;D��zM��YK�o�O�3�.3���ݛ=�����Su2����oN�M�&�j��{Y��n�</�I�$�+��#��gG�tC�k?1��벷7��l����r���_���Z$ʈ{`a��ؗ!��e%���%�Æ�T�J��kb��m�g��E�O��h�<�b��>xI�o�ٞ/�S
���W���i8}X�Rj_j2Pۆ*BVs�v�;Rm��i�h�Xi��.�*��L��1 r=�M�B�wX E��B�(����Npjǡ�gh6�y+��p��Q�@ Y9
ȚQo�5�4�b�
w#3N��Ɲ�n�@4-�u"G;GlG��L�����!J��AT���k/��A����3�q�0?@���eU�,���8|]��˾2'���:���O�YR/��� � �<PO���?�̕���([��i��ˡ%�3~P�{~|U�0��)�]�x�ൺ���Ka"�l:����������_� �B�2�0"�}�Wǂ%ٝ|��U�YJk��-%X ���x�[�B+�w)��d�)���ic>(8�º�%��^Wd�T�8k���`��5��`^Tòh��i1�:A�&0�)�#��:���qE�O2�7:��-�Cr^��~ݱ��Gy#1z�J�5+c�ă��b�W����������D�Z'��nץ��>��j�;!��]P�E�Z�2]!G늒Z�D%��^s�ҵ=)x��G��ꃍ��[�+lϵ��a6���=�8�̮�-y9����R�˂���!�z��h�n���A�G~������6%��;4��+���t�����8�f��; mY�D0�`p�+��oB#��S^�Y]�:�t��(r�]=E�Os�
|�>= l@�Ȗ��;�%;�Mmp_�#F���8H�L�gU�J�4:�а���Ĝ��5j(C�5=�>���m3]�?�A�����vS$�}ф��,��_����X��v�TI��'�7�����d����	��\�%ll���u�~�{�R�B�1cr/UnU=lb���-t7(2����W#.Ԡg�G����{��aIsc=Bl8y�24\��R]?6�.??��\F�v�9�ZG)����k�R�Xkf���݅����A��L�+Ot�R߭!�8�S4^`1��+%?Vj/���ڮ8�A$��jK����v0b;�Wpט�Z�(�Gg���0���F#7��)l�o|��R�.���0J3B���>��Fۀ��S� ����_N�E+8im�Bn=P��M�D�����Iw�Ue �/KL|�>:�VS^�B��9*�Nr�[�B\×���!k1U#Vry��~0�}�ނ�R�t]�D���7;�l�c˔�G�OΉv��8ɹP������c���ȵm����=��,����T\����9J<�J�w_����K��q� ��bY�/B��H��lo��X�D��H���g�p���x�{���ة��.0 ��9d���)dO����s���+��}�%�D��$�m�) %utۅO[��m�
B��J��|��
�F��w^[�t�;"��z��.��m��T�p�2��O�=X�ϰ?w������nw��5�ϟ��)�[3�<��D��NM2������^��j[��v]�C�U����/Q!��Yxub�G���p��R���X���O>ÚU3���i��ɨF\5.v����Ur��*]����@�*�3�EY�3V��I��.VK�n]�!�z��Fy�ة�켐���	o؇��.?ݠyO���x���g�4�H5��6a$՞�S`F��S9���W���<X�g�Q�]v�El21����^�I�vn�1oM.��g�O���lY��J4i�a��5�C�K�کT�t�h��́������O�l�O��A5 �#V�[qZe��3��$��9,�o�1�*��Sh�g��؆E�KN˦��i�&�m����v7�V#5�X���-ǥ�苝�~oW�na���7 Z�En���l���m`U�4�xf��j8ֈ9�wsXs�(aĵ��#���C����v�w@<�v�jB�N��ޛ��}�'7�z�+��&4�;��0�{C��>&�#m}����d_h&c�Ę4��_�_��W���}q��%��p8�|�K)��w�_+|�}p��*���8�[_�����Z���?��GTq����K��!�]� $�oRD%���q��m�
��#/&�>��#����zK�D�o�"-ؔ.��&�DA�|���UD�3�w�)B��Jͩ�Sd�2�o*p�����u���Ex)���`�������ѧ�@ū4"��~ز>`���ӳ����fE��ELmQ˨�������C�/97l��K�_jl	�JHp/[#�*���W}/[6.�L����i�$E�4K�M��t�������NM���J/~�p3�= ��q!���S���1j�Ҁ�3��73{�l&�ay�y�&���=x�P�;�r燠�׎ͥWV!��-�jw�7r��{����w$s�
9*m���/Ho{��r�Q���%ה���{�3����u@��/н��������k����Y��?:����A4���K�5*E��K��yҔ�B��]c�߿'$	��� ���;e�:��a�뉽����u�╀q%�ރ�+�nΕI�������v�v3���Xf�	o�����?��~RϺ��m�}�=��g�C@�3܅����u�����	M��W'��y2'<���l*��:��77��C��%���_o!au0�3;¥J�H{1�m���9G���sJ��^�F���eR$�x�{��u�$�;����+A;Ѻ��/0@�!AB��������L�o٢�	N��3?hY�OE����L����nD���k*�����- 1C��E�I��,�h���'�����D:"q��F
d�&ͩR,��>�Z@xN����퇥�:���������f�$�-\���@.7a�{C��݅29���������Gcm�ar,�k�R?��[ tz1v�[��agO$�Ҁ�Pm�Nڑrl�'G��ёt��ʐ����T��@d���loj];C��Ct ��A@ӭ�J:�����0�
\��.�������5�j��%�#�L宲���tF\���u�;��	�?�_Bx�!��E��u��ؓr�R}����j�s]l�m�"�ב)s�<j*�զ�>&1�^��q�n�<�=
�N��S96[�FׁWY�	֔/���ײ����������H�8�%~/�FU>�3ʎ�w�k��4/(�a/V��W���l�cS� �J��W����[��,��n���������e�''��*DŐ�kj�bC����Z8�l�,|?�����լ$-�0��Q�iy���N�Uӯ���8F��n|xE ��7��ʪ�	����0�lrѼÉ κ}�Q�)�U�p�������&���l9�����+�b����{��������r��6�v�� �|�8ʹ��c��J�ׄ��X_��g�ZqƤ�b�&OJ�fa�O��.�ˈP ��9 ��v�*��8�A�~~��-ܧA֏R4�0Qϯ��3�ǹrG��9�
���8��d�,=��a���1�Kg�dv�G��e������T�1��63ރ��u�з�+�A�B�˄�^n�e�)���s�4��kĆ�'Ae�0�����^j�1�.|�FR~�G�kID�A��a�����R0���Q�G>�m5�9\%r���x��&���p�v�B��ح��7��'���'��隻��זM.v�$��6����Psh�(B��uZNc�_Y�e#a���˒�HC���� E#B�kz�n�� ~��a33�P�,p�P� �k)ޝ��t)l�5����?������\��^�"����ЁF�i��J��(�/�V�F/lю�J�dI�|wK�"$��%h��$�`B�eS[n���$\&�]��`��0�1?`)5����[��nk�^�NP��IJqN���
�������J���!Q�����h�LF0�]g�}%p{��t�Sa��2"L	g�����s1k0��0�w����r���f��p�^`@�]'���S蝇�R����h`�@s�x�Ѷ\�/A���^_����ѳ���J��Z��e-�eJ��d��C�m�h��소�, i)�4��Ժ>�dUn��I���U�#̙S�Z'�.(���+ʹ�;&}]��,�t�[��ؘx�q�5w�6u�l!�	X�'�-�!�F#�B�S��h�~��}i2߳�A
y���2�=�*��״%M�Z�k���;;f�Yk�q�AZ~�ДУ������㕒O�p�[���b�<r����zrn�Ů��&��JP�xȵh�W���;j���mb^�2�L�簘��Ƃ @�E�Š�z�\�\R��~Ϗ�(� Ŗu�7�,�A��~R
��.�iկ8��+=�n�;~��&��4*��F�{�LLϯM}�����d��{��K����<�c�Y�1:�������GF���5q7�GU��$��V麨]����J�tw5i}�{k��5g���OA$��[(���'��9rN�ң��G["���p�����4���
�&�؎l�=��}�T�j�\�%?䐤w�<S:۬��$xV���
{��,��S����8�.p�"�0��G�D& �F�9)I��q����"b|�/n�s�f���2Ԥ�*\u'���#]�P��79�o��%���Yѻ|r�����W��΄ً;����̉�
z%� �S��I1I��Qbi/ꇷ�h.dC��;͞�wAicp2�-�<�B�20w^�
�k(�[�PN���R�M��d�$�����
>���Ө�?C�6խ���S?.�������L"�z��d�����vHp�u
�3���)a�8\K��H�`�H��Q�Ax�e1FAI��D��l#��f��J��~�[W��%$��GxWd���9~�LE:���_� <"��EX�U��k��y�q�4��3�`w:�@���c�9�A깡
R`�Եd���Υw�`�9�%sGSn<r��9���e�z]�)�,En�-��;��8��x���W��f��)���>�A�}ψ���@ѫu��A��O��nZn���d�f�Rw��%S��F�1�v�־��ɉ��6{.p�6�n?����i`�k�I���8�C?���T�1����%F�s���3X�[y|�4p`"�̢��oy������쑅�x�b�����k7=�Qh�5�ҟD=s��ίV�)��~���X��A9��J53�[Q��h,T�����%]����}Y�J�)�:%9D&��49�H^!��Pu����A2-���;�`�S�ƶ��Ak�WPž��ӱ�;���W-����$�YJCU~ �s�����\�����"����!�i9���-����I�R�3����I���, Q�����5d�Q�6'������M�Q�6�51�3�M�9�}�X�V
�t3����E���tk�л	�9;�E+��U`�n�������c���B�Q��)���~�o��SQ�pǁy�߅��Z ���&��0�=�yul��SRL�z?��n���K2���Ů@V��PB�`�v�4�3Q��zxjڟ���ƪN��&i"��Y��U�i8[>7�x�_���z4�W*�Ȕ�q3��	�7������w��^n��Y:�\q���º-�	
�4m��ӳ!y\�ֲ�a�+�W"���N5x�e�� �Lj��T�9�*��$��0��MP��F�I�u��#��C*�8a�~L0�{HFx�8���v�h>�X@d����qf�!�-�s��/�����7ld��	�3��?
tְ��ϳy�"�����pC�k�7ӷ�s���n��-������?Z�O_lG#����$��)�5Z�;�eH,�����ӏ�vjGߡ��)w8-����ʨW'�q����	>�SaJ��D�A1P|�o��p�
�_tH����N�{��P�/���w��JoX�M�챜.X)22t@^FS�Bk*�/f���G�HYw"E�YW��q�n��)=N�F�W�����#B�4N�MX�Ca��>���3r@D�]��)�V�8���b�ŜNu"g#����Z�^8�OI[^z��	:��'V�
�,Q�1}i��M�7��d�ᥖ�\g7��㚢l�L��aĆx�F���o��pA���[Զ��4��R�)!�Xh$�Ɠ�DဟF���q_���p<��]�h�w�������z�#BV'��tf�o|]m0W9
_"GݐN2E���+�0jkr<YI"{wZ`v�NT����L�Y�Vd$8O��� !���1������:����2�e��Ȉ�҄�2���M�_E4�E8|��xi��&�AC�B�z/��VL��JQQ)�����+_1��#�*:��P	�ێW���ҒEL֨���0>T3������˸Fv��F�!n [��eU���8�>w����1�k�pc�� ��X�{�����4	";��@T8o�wF�����k�����cp�P�`�pEflq��b�	N�\q�2{�b�]��xe����lf$��<�3=�7juC�OkzK�E�/H!iU���T�������ɕ�pl�O�j&�L� d��TǞ@�!ry]�쒏7M+_"n�'GN��F9͞$�^]؂��i�����4��,{nf�0Eϟ���^֜kV=�\y�i�'6dORC���'Ɯ�H����|��N8tNsW"Ú��='��T��u84�q�p���)�cp��vL�b���O�Tg ���K���P3ʌ����ﭛ�|���j,A�v#��<��zZ �:��n_ʬ�����l{�45�Bgt���t�W����D4�eD~H���3+@tv1����d��FEa���¡�ͥN��T���/��	*�h���X���4"n*ݞ���
<���g� 3��Yv�q"3j|�O�˄����M)B'g��S���"�^��cb����|�0�(�@���[��9Zʒ؃c���/�n��X�%}��ʕ�=dKԍ���&�Ӛ�͵�5+ڞIB!�h��[�/���`g�U�,5������܉PU[ƽj�T0�P�c��-�l՜ޮy5MA��ץ���y�����Bwj���Y����Ј�t��f�����*j�p�=G����j�#5� Uո�l��7�g3������	ڕj�k?J�$6�����U2l�R�1�ZM3/������(؜�)�1Hb���t&;U���-��y�)�Z	q` �u@�����v���m��P��׌>`���D#�������w��
X�������Ns_֩�`	����\`1�G����k'�]�v��FJ�$������7[�z�Z��s��ؾ�	�A���fX�-�d���ޗW��Kv$nX!����BDSi��P�h��솬��Z�@[�蒀�Eh��q�T�����vd��%	�C^�V��V�@�Jy"_��j�����M�`�p�4���o?5�7Մ6��H���|/�~��&_g�nKB�Z��qt�՝�E2d�������5����ё˹�U��B�Ai�sR���Jd��*E<}5
_H���&ܨ]�D_���g#[�.�8�naۼ�n7��Ợ�V:a�� S�Ol$��&11V,0���7�@�L�HI����A��#	UG�@��q�&��,���̥�oK��{Y��Q+� O[Q>2�?��#��(�?y�����YW�hu(� ���f�Ў�b.�~�^4���h�R�`	iR⁨�A_���F�6�xK�֓���dR�ɯ):_qD>h|�����q|Gr��D/��j��j��$ɣ���J|��mI+��
���v���,47H��0�[� 2����GSl[���+�GV$�,�t�	��=Ou��:k�P�]�O�ձ�X$^w`�6ےw���:K4Μ�}�+����G���,��b,-M�mu,nu�n��n�FP\05��������d4�z4��ދ���v�a�/����5�.Sx����ҽ��!�յ����D��P���P��S24N�A<ߟe�����Aap��� 7l�QS�n��]GEő�GȄ�L���a>p�/��C�h<<�HN��y���_�qD�o�-i4��,Pi���C{V���W��?�/ឯܒj��(��Z�h*o�O�O��c�$�^�=���*�9�����E2��zIM��7_�2�������TͰ��2,6��j���	��RC�F�O��m��t���L��>�o5�����?�Fɼrs!�*&��.�}�s�ے��P�iqf�ݜ��]�X�We�Z�0���n�*��"E61z��1�*f��~8��iP�fz��g���N���8?��Ųd�[��UJ>̗ x%q�Ӵ�|��sN�ͯ��wf�Z�c"�U������Ҡ<��
��b<�h�=+dfK%X& �&�F��	,�H���X�cf��$�U�O	Kl���Id�
T�u.W���h����/n���+{�hj��id����D�2�?gy9�lr�2)W&�D�e��R���a2��'�fp֍��4#�����3gu��K��{v,0FK�����=��^�H]�61�8"�1j�9��"�+��P�.�9�y9�*����غ�\����t"s��{'�%��l��%Ƃ��w�I���|5���ޏ��0Lk�Q�1�nKl�:�)��$�����	�w����MM���f�c���aȶ�*Hig�a� �%e�gEH�>���8Y�f���	E̛&��ɽJn7��ONں�-��Kj,�$���8� �\H��ДaK����.�?��0Gk��,�h���6�\�.ϩ'Ϩ�V��&������.�A.��M��H]}�(Ъ�o����`)Ġ��7(���w�)��� �}���g8���qh�Ԃ=>U�Oc���<kRw��֪�nK*��:��ط��C�#�����e���pKHEÙ�I�he����,nŧ��y��*A?/d�D�F:�-�Nu���~~��3��4������kt���'�D4x�2)�5�,�/X��h�*+�?�&u�8)�C����S6����qud{2W�	���	M�]�^���y��7Rkd{3�.m�57���Oh���o�;Q�ˡ���0ĞA�A����	�}b�m�E��kB�nG���NZ��8��KܡK�(�+��yG����ۺ`����8�.j�v~/�P��H��0^4ں^�����>����>X!����g�@�ṳ gj���|�ƚ��I4�2jg��2��9�8��%���9T�>�a::N�8"�Ao��<���o�m��y8�0�6f�-��Z[s	�܈,�w��|W��k�"��d�ͧWZ?}���l��G#�9�Y*oϗ鉢��in�B�x�s�d���j����V�1��zP�9��Zm��i�{�dr�8�l8Exҭ�O�8#��2������
dJ��}��`���֫F�T"� �ɢK�X!o3*���o��N��W����֪��y�4��y�'�;��k�Y�l�v��*4ABsQ�P���/f6(��ۅ� ��6E����L}P�j��K7�*o���Hha`q@�]!�yf[�ٴq>lKn�'XчZ�;=�^��i�����2\CW���v�N�L3,$ϐ
�oedy�z�e�y�����U5,@c��g�[֊�ǟ��t~2;x�ҢR*�Z=5��F�!]u��up(v@��ͨܞR{[��V
x9��#��>��+��	��~�����U�W&��1�ʐ�\�o2 �.�l�����¶�]а)��zɳ��l�����҆�R���*?��]�L�������z�K�������,�����-nփ+�~�0�A@q�Z;P^ƄR-`�+O�v���	n^����7�ÂBI�҉��o? #<�0��j��_a�B�\+s��<,���kK9O�
�I#��U[(4F\�����JHdlf�Zc�{ZqN�����]���v�'�e��>/�ۯ&}�E>Se��,���n;�'ϸ�L�`.�+.���D|L�T��hEe��EU~W�D`����6��
�fyG�G�[˽��G'�R��67��;䖎��\��pe)���������>�go�Z��O�]V�2���tkSxeٛ�:����	������8��x���(��З�c��kv���I&��A`K+)�i����:T����fa�MP�d���!Z�O5�f����F���M�LW%~r�.��|@k'��?R�=*ɿ�WZp��O(�S �\ՠp��@tj\H�2��9��#�+�+s�}77���!��\��h��&����Y[�4���$Di�y�#ҫR:�\yc���8������#Ӵ���K��n\7�*����%��_Ru�Q�U���o��[t.���-0O����c#����~\�O�1ŝ;'F����3�"Ľ���+��$:����'( ڗ��M5�����PU� E.�D# »6���ͪh`{��_e�����">Zi�7T� �@������~}�p����ptX:�/�x��Ծ��CM��Ћ5�׮��WY+j�bw�(�e�rI�f�h�o���
�WG��.�*������sz䷡TꔾМ'����2�{�Z�o�<DD�!�+z֦�)�.С����_ћl!��EEbT�]�(��Z*CFux�����Dۃ�3h�Q4�����'K�<s-���dzUg� �	�VuQ�L�r�NF��+�����MDў��V�e7.Po��؞UP���P첤�J|��o}�tVt�x_��'�ܞ���1��Bҧ����hg�2 z�K]On���&�Dp�N%�%ȫ�����L���Rul�P�
9}p}x�r�[Ɇp�9Ss0�1=e��[,�Ǘ�`�m��Q+G[���9R��-�p"��y���>"כj)�)�zA�;ʖ�I7�����z��3�{�EUP�K
@�����-���U����iX D�-���b�NfGaN;ƻ^f�u@TV8�z=Kq:�[�Q;��b�͋�o~�����w�����8,tXQ5:k�е�keh���p�/�gc��8�x�c/f�M���	邘�v{�3�m�.~��`<~b>�GH��49{I@��A�v���ٿ<��_B����T�����+8���Q\���=U 7����%��)��j�L��zP��m����g�������xQ,ss���7�4S�OV{PM&X�t�PQ��a����w:[/��Ы�S�<��l���w�>����9����I�y���i<�GK� =Kݶ�H�s1��\�����T��3U��/�����YQ���Ov�jxF��`���Ɗ &��)�P�E�|�"0�V.d�� �8�x������H�h�SdYLJQr��^9��^��Y�h�w^�zG��l�@�w��Ev��*q�� wjɞ}�����:{�v�h%���?S��Y㊏o�-�)v���]��᐀AD���-3�v\l.3x�ϸ&��ׄv	DY5�����핲���(�"]Șn_�/o�6�閚�ť/�L�9��_��ϡ �) �G������y ڱ}�r�W(��sE�t�IO���,W��0�1J����8�\��B]>���}�g��i6�ƨ@�a�8�db�v�F���t�5��0 i�[�.꽰���X}/��D�ч����G���M�}�"����7�hD��g㉯�D�2!s�D+mk2�"~��F��=�&N������;X�)�Ǩ���r���"ָ,��ך��b8�l���*�Zg=�崭���9S���#� �F7ō"�~�LMA O�u��ɛ��RB�U!�.%ϓ=<���Wzt�����x�(���zXg�Ϥ~�����/k��u�bv��~�l�R�'@ G���#��"�N�I�	�X=��z���y[BSr[�̺�V'i��$eҦ��IU�=z��N��
t�Kѯ�#�e�<�i�֝����/�1�58�=-چ��?;� r�l���R��=a�>+�2��)�d�6$�f(�7��Jz�\&���󇙅��W�.w%P���[��
D��X��/'E&!��e-�\�9r�.4������ɢ�%�պ��jK�լ�����`�<
J�n�'42�' �
���"Rlk�>C85�ˤn��P�Dv�oZU��3�`[�}���ܘ���:Շ�M��	%�����F��s8�FP���>W�(B<�I�g���p5^0��_�p��]c|�f�k�~��&/h=�]%�U��
]��t� �x�b�n�«*ӟN�3l�x�O�5��7��k�9�CЪ�ƻ�7a�dq�#%�֗?+V�J�"�ʿ)p��5��{���w��Gz�N��)�S�3���x��5�+P���X��sB,e����!\��g-����
�ɔm�v������L�F2ct@c�6�G�c�	/r���/Y�^��ͩ�sϏ�gZM�?ɖ�xl�{�0�"�0���|<d��B����c���cYv�w�+�F�SH���q>�H K��9�
aR9���O�[��2{K��(C��b"�k��cԣt� 8�h{Aځ�Y���*�ߍE~��2^k~=p��5��	.mt	燀"_���tI�q���Y����so�0p��~�᱒$cSE�U"1;�n��A|p$,aS����������f�t�����Wk͖���_���e�����j]�Wy�-S:�/�ES&�@���pUˤ�e��~
�Hx�]�G̉9@{�C�Q0%��y��FE����s˪�Bs�$S�p�\b���F��0�*xm���qh���̋@��~f��诛�/8��G�j��3#q��,@�K��ɸq%lB㿺��ꓼ� ����pl�+����]�x�}uӁ�'��_z�\��ן�"Y$ڜCQ%ٳ���(����4�9(#c/-�Kz�4~��sS;���r �.�Q�&��y �L.�o�u���}	�&p��(���!���� �����������`8��"�!�y|Pk�&E���e�_�+��"����C�~����iq���:m
����ԅZ�Pm^
��G�@>���A���PT/�9�9�
J#���儻2��l�G���!T�����<29Ȳ�o��?�M%��AǺ�w���nI@��#C��%�Mp�3_�S.��, ������h�����z�f��w��K��,��4c�q>��*=�}A���!���Ǹ��5 #��,�O-|_�����`�|3M��3=auY�/PlJ����9�*�W D�Y|��_�R(���Ab�ҋ��`�D��3/�0`n2���0 v{�QF��II���p�(��Qi�yݐJE"�Xs��\����#T�)PZˤ-�+�~۬&�v�q\o��69ʉ��ն6bXs� ��������`X�$D�&p�r?A� �̒P=��K�7�l ��}�8OQ<jc�y�
?jk�j���0���`z)��������4O�����C0��*�F�e�/�N57u﵇�y���z��7�"]i��>���rX��'V���%h��B���D@d��j8���{�2��[Y5�0�����]/kJtX�΂$i��g �RE]�J�d���,��mg�Ġ�ݡ۞Ɩ�P�i���,��, HeZEP��Q��~új�s�6��T�՝c'Q�S:��X�t�Ye��=������RA��l	�2�O�gl�p8��s�ȀT8��O,�-}G�W%T�P�M�t3�&�����v���T$��zS�S얌1BL�6�:�%��x������B=��yR��r��E�¦[)��81{X�w�{@$�B6Z��$s�`�Q��v\��OU"��yO$M�kX�ઑ�IbU�WELE�f8�����8<��<b-K����ր��[]���5KFi���]'�Rp��?��f�N�� �?�ӥ�P]�=����n	Êj;��s�V��U����=ǩݓ�k'��C
��	�N��wef7�g���a)�������u�x	�ػO�ɪ"6�@�XRHv��f>%���j
�e3�v���v������i� ��Le�GASb
�ߵ��'Qq�?P2�T.hAR�{��K;�����:���ߎ�.fѕRp���!��t%�
;k�1�ŏ�z |��^��#$�G���k@��r�t�,)ߠ�R��C�Z��*�ew&�J��\1$f�j�)��+9""$�#�_���m�"�c%ӯ>�(϶w��7v���@���/����&��[�}�d�jG_����5�>������NP�H��w�d�ș�k����P�i�H��)��Cd��ة�h�D�����!?�EW-&-<�m��B=q��1��B#q��c�}������,�f��ϑYFm|���K;��2��U��(@��*u�w � o�=:�ӽ��x������h���V �mW�,��ҹqL��қ�wޝq c�ӔY�zc�FI~��0�Z]R�0�.�	:��+�ř��Yo�%8evT9�]���+�C���������BQ]3
�/�bf;ų��K>(��3;P����B�\���\�Ҟ>5�F�l�.�\�M�����M�fBIʧ�%A�mx��p
X�o[��'�� �d`2\��	v2SG�����dcx҆�㋢2�H�L��C��ݬ$E����X���Y�?�]���F���aF:'��Vf�P�B�h�U��b;�*5�%%�8�&�K�S>�g#Hra+���r �*�,��|�]`��W��#ɱ�Kx*����W��"��z���Ot��#f�T�x�,7�7�お�T�a��,پ��ykGC�V�m+�;$�����J
���W�-����#��t�^��y�I?���i�;�{:�sv�Nݣc���<bt6կ�Ȳ-�Lz+HO�/j\'���Ct�U��5cxOO	9r�I��cvb �!c�E>��,��n�L|�4Z�F;��ǔRq���l�K�L�wfG�	���y'd�ʤ���>�M} p�����Zm2S���	����Q?�I�-������'��%)����x��h����(���ʁ��J6?QF �}9�7��4��f�@?�{
>��P�=���/�e�9�E�WL�S\ Ϟl����?��L��i�8n�&9-U��N�u%�.p���Ҝ$��
=;U��o\�Ͻ���[_㚩�� �t��jhE�49Q��	Ŵ�=O�k*e�`�}c/�$��@B+�/�*ȿ�0�Q�a������rմ��*�	%���iv��l�\'�BB�&קcmx�䤨�z�iˍ���*+���u��S�L:�� ^�s��c�΀@�Ϥ�oK0aښ�PS�"0s�N�buީ]��Q,V��>��61I�έ@J��25��Ǐ�)�x�'�$ ��ʜ��X�������DP#>�{�R&��*�x(�&t�å�[a�Â;�D������gO�!�R����C�x�.�?$*q��������ߤ����XK�X����<v~��u�=��B4�cI��c�Ic1̝V7�G�r�� �\#vi��G��N�NU	H՛� I5�}��I�Vs�й>�2��{�]l�図A��G��_�Zk��c�u��i�('_�?�s�GH���e��E�C�T)�NB*�0W�{�<z19�F��2(\�����>ׯIb|6z`#
�t�T�w�Ri�����[�U�3��&A:��kVzEH�HpͿU��q�9� >�?�nF@��)~�l}���g��'�[�̑�����i���V��+��?����=�苁)�%��|���k) �[�q"w�4���)j$�QXf�;��S�x�E)�a�Ω��z�!�5���$#OD[�g�X[����	=�G;t��p�m.&2�	��<�Lb�����Y�w�B�/�R�׏�2i������{�x�Oh*�����Ջ�K�}���'�����f��B�Au\�cbl���.���,U{ڴ�<�"d�w�X����n�]B�]-)���*�Do��-����nnyD�>T����a?�[S$$c<�f�,a�l�<���i��VY7gy����  ~,H�O�6F�S>�(�fN��ek�B���A]p�T&�:Z'�
a�W�w�'1�q�B�V#ɂ�
3I��ϬJY�0!��K~�[%.��(�f�,�_��덆���%K�n5�M�D��hږ�ק�l�/>T�'$%&-����� qy��:��e0X�V�v7�_5�*	�zb��A�!��ٳy"��Z��C;���4Lʐ�90iK�4F���&hΠ����1��`��Y���Ц�{)��2c`��uN�B�f�P�V��R��j���7���9��Do�P��l94���!�G�%s�I���c�������ߣ]y��,5ez�m�K;S�v�Hee򃺀pܒ�H3AOJ��(���ՙy������d��w�}+�KÔd�\]������~�x�Y�������6�ҝ�=Ï�!x/2�<��0������#I{��U�|X�z��Vm|�ҍ��Z�1@�����?�7?f�Bμz3i�.?���Q�pa��+?�4���
-X��$%H��).D��Ỹ;���\�_;�&��ʕ[<�S�����x�|r
�9D�s7h<j`#�Ӻ�Plhe:y0.r�l4 �T���~�Y���@6�p=�٦�-wE�d�R���	�q�tP�X\m��ԯ��8m�!���� �^������?���Z�<y��*�|� �i�f^������t�͙攔�:!����x��4c0��Id"D�#���X�N�'$8�6Ƽ�/~�5C�V�0�w��{o�����$���|�f��gV��-�s��L �pG�ޛc�0�~,��In�z�\ra'%$=���CLV&
O��2׾UX����� ^��<����1N;���\5�f�{��h�E������H޺�b6vq�\��g��+us���\P�T�|��34�7z���Cp�W���̴�� dV�@�>sH��i\4�j�	^�y�����F<�?�^-��5���5Ȳ����F� �4/��rޝ+���)3�*�k������(5��	�e!wKR�H�	�9PS��C� W]V j�4���^i���,[y9?�;wX�4Q�Y��-���,�K& ����,s���A[Hh�n��໅\됇n���4tP��^��Ƣ�5#J����7R�*m+��	�0
CԸ����~����I���X�f�s(Su��+�&�2 ���(��d�@<�EfV	O�n!USu��ޞ���֊�J*�QxU*\����=��^�c���;=�����Z� ��c �p=
�#�lkp̍.�p�AFҚ(�y,��ʉI=���p���3maϧ��q]��W����.`�\�Ŵ�9{J~�o�1˚/QhŦF}����m�d6�舍
����a�D����ň�"f'���Rb�i2H@�*�T�=A�p���Ww�S���!`e(����0K�S���������B�]���'R
��C���xb�s�Mx54.h ���X�e���d��^�˅O�<�ԋ��G��Z'0��d�:�(c!�U�҉��O����,�JH��~�^٠_a������	���Ůz��:4?���y��Sd�ٹx�wgJb�ɤLڍk��i:��R���D2�AN���v
6�eS�ݯA���7��6<�;%`\��;��k�� {��� w�$E��ôދ:�s�Q\z/��'��v��!�\
�֖��D��G$�[��
�}Kr^�xu�$�	^���. T��;��3�?#�I�Q��tK�X�o9����~�{���W˘=��YR&s�Z�����nfپ��ϭ�@����D��~�*a��-�5�I�hx9yn�+�jZ�ި ��iF`ف��e��$a���Q˳��(��:V&X��W<0�<���:��? �8�q���|��w$����r�{bp�MS�{)�j�S�	h=�<�D�% =ɬ$��Y��.�K�.]�0��m��o�]֍��$J���c��TOqT�:�Mj�KIZ����Ĝ��[��&Ę�<{��w�u�3���O'
ޝ����������t�=�(곿�̬tѡ[��@q�Փ��T�v�x��u���D�����Ĝ��]
�G��� �k�	�w���T ��]
2�IҴb,X���=��5V8��NO��9��~Hr��!BP-�c[!�>�cn����$C���By�u��YOrn�\h!v��`-�6�kEFd�)H�����Ƞ�=4�K�>��6�RM�6���LZ��J2Eх�IK�hڠ���(��@B�1�_��:Y�"ɥ��'�"�N�����N�����-���]���!�yL�#�P��?�h:��D�ά�J��02������k1Э�0�I��R3��x/�r/�m/��өhS���_�˛ե_'6{��1?���v@տ)�l#ji�f�2��^��>�4b!펺��!�K�����|dj�uM�������?"�(BO�]d �Ʌ�ݭ	%�4�t(�x~��ruJ
($��3�ݠ���N������k��\g��Xq�uQ���2nT��Ĵ�4���u�+�H�J�@���q��7�_�F���,�-�[{w���Ɖ{�
a�O]�y7;#�v}�>�^�A��yl�v���m�,?���U=H5HdG�DCO�]�~#~�ֽ���Y�1�_Y75��e`W>�TK[x!!�=Z�%�l�@d��>Dti���F�#�zITa���;��U��D���#r^���@�a�.�*�@�_r��#��`�k��0�M�c-���nY�%敖�+8H@�4
�Pf�S��(�*�>`fir��G���v�Y�BHǘ���#�T�+R%�g%�GB�7�Pc�E���B��y����*%�Y�@��Q=�gK'�ױN����:��*D��݌Ca�:�3R/�%��-�ڜ��AeΕl�v�NҘ��"�8�n���@��Rޤ-J��l	�v�|�Y̙�i�%@y W�(�$/A0�����]�?|�iv�FLdCɶ���c�l�]u��!�Pb�g��|L��͑j�J�{������T�뎂t����T%�X�*�?x��t,�kb��POÔ�0�B�޻�PY���'ђ�\w�����ѷƧ�A7�V���o�zZO,��;L#���2*�Iq2��J���Db.��(����<$�c��YP��8VM��������/Ɉ�CI�o����#���Y�0}�e�cǮi����l��Q���%ŵH֢��v�c��F��ZQB~.�
E�Bu��&h���DF-����i�-B�(��G�%(��PP<�[[�?��W�*�tv}�F�T^{�]@!����A��$���m��2�A�sUex�����q�Av/�{�E�h�H�|uiW2O�:�����j�cst�⇣.��~D'y9 �,���]����X��91)x�ޖQ�q����G�ܪ��9��f;���N0D$��=f� A��8�>��Ip�SR������ 1p��/r��p��P�5��y�*�ċ�D
��ԇ�.��9Ǧ4v�%�����8��0��՛�����iA���6R�i�I ƴ����e�`�C��j�����%��z^8-��P>����/��-����f��;~���*�I"~��(�U�����=&�T�R��}Y��!�%&4�U%�i'���j4=hIq�g���i�����mѦ�l�i���e�XQ�9U�<,���4z�Nְ���2���$S�n�_�4�c���i�� ��@�b�d�"���� U��H��&Ia��Jy����b㸳����������T[F��yy&�W�C�6�Q>\�4fIM9�yWmt�=*��p���EG�%�r8���K�N]�Dv���� z�
(�+D7=�����ffGJ06,s��f�%�K���hp&�c�q"�MI��t�5=Mp�#Q�����c0�gaA,����K��Bd�Z.,ĈY����n l�
-a�>D�kS�$���kE�MϘ�p��8w@/ w�L���S9�#y���=�sC97K��r$�ț���;v�v��9�V7���tH�S�U�"�h�)D�&�_�9&QӐ��E�(�y�m�1��ۚ)�Ҵ�H�Su����d�^Ӱ�e��T&�|��u�Z��0��q����|%���{/f��U�����\�2'���s۹ǈ�}F�*��Y�՘[�YL���Hjw���!Z�����:�նr  �<MI���\A��[�����kE�����n`t,aY��[�D��2� ��F-
6�rdu̦*��h��.��Ja4�+�y��q�<D:"����q���[j�=&���VA��h��].g���fN`e�4�K%�S��ŗ0upN�X����jQ�]-��6{��C%6�����a�����K-%�A���ӵ����[�k#��f��7(�Nܛ�,U���VV(�-��p,�(��GS��C�I����?�S���$�"=
�<�ы)�׏�g���=�<����ɋ�����0p��6��U%��!����]�*&"�7�
��2ǰS3��Ғ����1��u�c_��ۄ��*0E฻c�i� �ۘ�����b����7���A���-|���n7��� �}J���d@��s���ܧK��V��Y�v�!冐3���{��~5М��/�V.97 �F__)�8�Go��A�U-K�M)\1��Y�06����ܪ�Q_.�X�S`+J*0y1�\H7���ix@	ע�<���$�഻�F���'@^�U�r$�r���
 #�U�;��n�OD?O&�xS�GN�&)1��-`U�����f,��֍;�D��S��g�l�FKA87�$��Ez߉��`W��h�S��,n~re��sC�Rv�(Q���v��eL���2�A	���S�	��G8u^����xv3��E�`n>Wa3���}�HLy�k�UA����KH0G&��S��v��Z����4�W��`��!�<0��ڮN��}ȜP�����o<=~����X|���֥m���׃�dB<�Cw��Т�VP�:�ؑ#6G��|:��>�p9J{���g��.��hKZkx��"���<���ұ��;?f[=妢Zj����!���|���N�O/���[̙��#c^�����&"*��O'��n ���IX��Y�L�[C�|��,e/�c*�)S��%}"M����(�F�<�IТb>@��[/ &���NODw٭	�'�L���=i��Ă#h�A ��ۗf���@���}`��ӎ���)X�f!D-�>'˼���y[Ϲd���lI�uDID��y^�s�0�9&f�II'���b�Q�/�R��پ�5�T?��0$+g�b�*P�����O!�Љ����%\���u���Z_���|�mU�p�N 	,Sd�\!���׈�$ڌ�0�_
�q�|﹦��f�����A��(#!STۛ�EF�vD��%���3�����c{�>mkA�s�Y�-m�S��,RA�U����b���ʅ��K���7���p��x�w�*�^Z�a�H��w6c�W�4��l dZd���o���j��LAۂME|lK~r������l�N��6��6��ǶJ='�r�pF��F�+Bc����~��+�=ݨ�]A1GG6X6�`t��3���/e�����dͦZS�2�0�ۈ�ְ:mȗ�0���mDnf�E���ƅ�4=dCG��X�N@�!�v7�7��N����h�d�r髍zQ,��i��əq?��V?'+���Ch��}@!C.�`�oͰ��e������w��vH����陇IW��	��2������۹L���<No�:0W{�z.�()V������ <�K��D�ޓ�2��L��=�y@8�$��;��[���_�gc��q�~�1i��F�ϹN#m��^o���H��	��e����}^�k�4EI�]���MV��wƟJ	��Gel/��>@�c��?ԐaOzò�\�AT���+rT���O���bB(B������ j(7|N��v�W��x�m�d�V�U-�Zf������|T�xNԵ��o�<
�3T���tS?S&c��L#�d�4m~���
[�P)Q���@��i�U��)�L���O�wTC�7?�B
j�c��ԤL�f�Q|�u�N}�����ش�ֶ��Caœjs�\��a-�`._P���k$A�^A�u�Q�l�~/��h��� f����	O�t��DV�q^�Pq�9��@e���w�U��oސ��!�B��k��b�q%�qI���_ C���龫rZ�	���Єe�/��@��o@+M���j�l1{��݌�����&*�dX�v��9��ea�1�0�n��;H�P��a寴�`�j295?w4{T��\h�z�K=�2��-�[�� $"�l����R0����kU��H�H�uru_W��9i,�ɯ�~�pHrUN[� $4�Kr�]e����1���f��0�Y�#8	�r���z%��:�Ń��3^H�%����U�;f�({��>@��Ork��?i�#m�*p�T.�9�q���L�u�|ߩ�Y���v������$Tz���aYl��M�"m�Y�g]1�\x�`,sdf?�It��l4ONU��d��2�pǦ�O�Ֆ�A��ˀ��"�@���&ISڀ��Gk�8d���V�9V�~�k��"Xc:0����6ab;:Q�6��g1ܩ��|����j�zodX[�}�8@��Nn�,l�=t&�)��M��j���$�c����l�#�[�]*�7q#!�hY�S��pm�hK��Я�$����/�-�g,�]�vY��I��ʝ�x�Wr�:n��a'���
7ǥ����-�/�w���)|�����>���y8$��1Lr\g�o����O䩥y����C� 1�m�����|�I	$Q_D	�F�3�g*���#�@�;ͨo���ci[����������ޅ ���	 !#�e�$K�m�( V����s�(���Ke���f�&�i��sB�rr�j
n٤��<C�%��c�J)�L^�3Z)�!@{�7O����s���.4gm�L����6�檚����U�C�l�Ad��eC��A�QX�*.a�_��ŷ�K��3iZ�\(�#X�\q��B��j5f� ��a��:c/S�^�%2���]L&άs������v��[�S`y���R��+0��.J�S1��U�U��o�k��������0"�l����nA����W�#`�2Hje���t��,y��7�Ml��u�����ŧ��
��R�!��Y�W�ܚ�gG Y�O%S�Xv���,{[������������������ ��4�<�n^�;0���k�b�	�B�K��|3 ���bC��\��~j ���YO�R4@R]�������Q�(a�Wj�͘��Zx6�x��k�c�v�W��3��1����v�PGb::�6G�yzĈ:K�n>�ꁆ�a���5W�D��ޮ5�(�C+��[,*b���_ �w�.�y�i�[��s{�5o���ڸ��}�������8 �4��D�T�:47�����\7�\O��h��?�s��1O�R@S��[�Χ;+���lЃ!�`U��ӌ�}:an�n: K���`b,���X�����J��(�3�p��8u@�2Ir���<�r��]���R�/�;,߽��_�HȰM�lݍ�za��l�:�;Qi�ل�oO�����?���ȣ�D.�����ST�x���">�(�w�m�O�i�E/{��fO�0�����`;o�E�!�IT��ߩ8�}W���~������*W"{���E��w5������Tm�F ����3�T)���4�L�q҉�2�D��  �})�iEcc��ÕAe��F�x��e-Ԏ���2�܎���t���@^3�NG�����ǐ-��nV�o)��~�TD��V��j���ZŌ�9�n�:���Pо<u�IDk�(��d�a:�
,I�W�!�L�[/��&��f���P$�	�
��[d�m �'h��zs�sLU�<1*q��mcM��������H�-�dkT}��$
��OaI}�ω�s�sX��U�\)=3A����ٍ�x�G���i��8�B�؋���b]k2�����K�ˋ�\_���Y�J]�(� 7c+�%p1w�)҂64�Ǹ�1tm�D`��9��c)=b"�����pU�R�	���]� �3)�`IOQ"Z=RdHLE�U'K������fױ��Z�?�7Wi!�#57���U����>��F��6İ{|�\#�S-��2J%4�L��z?���~����� �H��^�F�c|8����2��>g����y�d;����f=a@Q�V0��6�	��<%��ؤ�=����Ή��_�HK��9��!o�����WZ�-}��C�P���#1�����r���5���j�ޟ��s�*h���x����z"�����s_�y��
���9�m��)��;��HyvjaM�#��,��c	�m�xb�i�
�l�FX�<�QS\2��3�,k��8�'�q�P�dv�a���ֻsv�.*�)�Þ�� �X�a��!����A�������ط�E?t˰N�52���[cl\�Գ.��h&<���=����A��\��l�Ǿǰ�����سfqr� ܔtx'au���}6n�3���$taa+�#(�΢��y- �X!z�G���,!~�l� �I�!��A�K�2$�բ��zy`�����_L�O�\"�
ஒ�L�e��g���y���x�����Đ���*�Pe"O�����L�<��<��Tc��¹����Vq7r�I6��������!�b��)���K�E[�h�]���?�6c��~S㘃|�h�]�?��m�9����y�"ű1B�K��� L�D�I`Z�Z�8C���y��t�r0��Ƥ(�FT��tx�iF���Mɍ���b`i�p+���J�D�h`�ȡ��0@�Y1J�G
�?�(�Rq�#c��;B������ �����jQ�Q���u���c8�e}{B���8&�8��������U��d�x4��i��'��0�T /���)-ݍ
n��Mi�S�UMčW�`�^@՛�!��Š��w9-���|a��F�e���M����fR̨��L��!���AG���ʩ��V�"�@7ʛ��z���7;sc�4�^����Jq��W�tT����n����Z7lkBp���K�
Jn�b��Y@#��f�I��\�愣��Gy(T)ozi��@��bE�_T۩��y��<2��F�U"�`D���L�ķ�	���'�v�.��.�G�'ޔ Uc�.�6r�ߗ�"�#`���6��GQ������	ǫFΛ4�	17K樚!�*�(�W�c�R���1� L�R;皣T�_ˣ��V��� ��RUpSO���b��Hl(�^C��fk�5DWPpvƅ8��2��h=6���C7U*g�@������7�O�&��+��G���䒰b�����k$�HN@.�L�q5�Q!�W�Np�k�>���6@�i���8��wM��Z��bm[��y�#B�Z6`Mxw���ѥ���;~U Ӝ-���QqT�9�ݾJ��,!A���`ݒ��I��T�'�v���9�Z��)��>�{����v��@�S�`��߬�x�2��67wڮy쵂��Y�[���J�I�[:s��U�P޴v�](2c>��+[�s�K���K��+)�����G����ٵ��OL�C�Ƃ�S�����b�j����b����b�:uSw�a�򧕹�1�4`oƬh���_�Z�w}@$��z�pa�<��8�GKR�hn�L	h��d����+h������4�|��E��_zP��K�!u MԠό�x>ߥSw���SQ��"<�)k�wV�][n61EE�?�K\� �m�*`9�<�X����!܁�k�`aDMJ����\�2B�"�X��0�!B��N��#v��6��a_M& �:VURp�&����Y�0.?6DPi�T�U�ౡpC:ͥ�%!��B5�� ܓ�6%{���
8K,xUq8#w�ЕN�>��d�v�AN�?��L�p���Y��Ha��$䡈8͟�Mo+.FU9.�Aj�� ߚ}��K���EF?|�IQf5�-wD��|n�
�0��`&������އ�3�1�$��;�A"Q
�#���z�NQ\������q/�i�I�6� �AC�l�,��Ϝ�p)q������[�͸i3�E�e�ģ��z�*`�����wH�Y�S���cYL�������G�6%��JS'�yd@3��?��"��2x�r�!���6<��$���z�������:�Y<KZ�3�ŉ�n�y,<Ũ/�r�����{FXO�8�uO�9F�MO����b�Kȟ���n�����E�@�E���9z3��A�C�t�X���0�	��J�+��$���F���}�c����Tb.Y�1�֣E/1�\Q��9_�ҘJp�����@&`��/L�!��cD7F8)����\�,�`Q?,�@�F���]�ԁw���;.�C�G{����2cn�v��`3ګ��
��mD?ǫ+�շs�\p��By��G)8��V���x��!7��Z1�8�����lBB�~��|�	�!r-�Y�Q�Q�񡏫���O�!CK������d/F��|ʽ��.6M����ߚɊ۹��5��>.(�ݬ��A6U����J������Eޡy�uz_&^m�Noe��hcY��A���J��u儁Ց��#�>��^�C���k��:��GXY��U"v=��Q���VK�52��٦�a�R�-��qD��0�5w��z꣕�
�#=���.7�����Vz���rq�H��O�HJ�5Ro����-!��1�U����-l��m|5�W�Q�5��IӸ�Y���C�&�4�����r@�2!����	>(l�9�&�(�$���I�8Ƞ��9�^ס:��T���n8�&F>Ǳ�9�߼�ӆ�J���n+F�:�����I;��e��mx�^�俽7,cj��FqU�M����OȲٙ�[�(�$vf�&��e7'/��d���?ڙu0���\`���NF�i�b�O�֋�W}�eӾ��C��MJ���=/BE?�\�ߐ9)5�5�l�����=���s��bj$@yî��z\i�y��.z�]���f ���ڏ-��ȃ�I�b;4s�,|��ݸ<�ʑ���A>��]�PKL�8�;�ċmV��+"F"X2ܹ7�xM-)d�����3�]�����g{K{�dX�z�|�����=����o���֙���r"�#�c?�5��c+��'fC��%�Oc?���\%P����m�V����)�A�P�ov��5h�Űc�"�+��Қ��D�N�X��F�(�������].ޘl��<��.��m^r�!�5�sa��T�����;
x�b:\u6�=	�hӡ��Qɪ&�<���&��y�0�+�LUzE#�� �iL��ncn���3Վ�v`�α��1��T�
�.3d�Gj�J��/CU����$)L�xr�n�hN�/`�DM\v�V�/���6��!r.鷌���z��4�0G'{��f���KG�o���[�c�f�쎣��}�P�yg�.X]Z��Uf!7�`:�q�N����D���*� s�*�Z��i�d��.��2�i2�f 2!��z�S���eْ��y�#�ߞQ恒�N�)����	ׅ�\�
�>V�turk3WG��]� A�t�W��m"���z ��J�B녬��l��>N� %K���	G�jYQ9oBɀ�m��i<�r�M[灟q��J��[5���"��y�3�b��D,�>�*�0�h���A���(n��Q��k�K��F����0�*� g�7?c�����D7HR��La>�z'Q���q�c{��~�	�,����EFC�Յ���$�KZˋ���_�65I�,��� ��m�����c�B�X��%8gM�u���&���߄��s��%'w���b��IV��p�L���GХ�,���0g!da�E�� ��y�����Z�,^��4�:M/�$0�
�����2�.�D� >�.�`�E�d�K�1���'��ܹ�\�b���� ��6e˕��y$���&y��^5-���@D��yz)f�X�c~A2K!P����M��1s����$���YaL���|9N~]MsM�ꞙ��H5^��(���w� 6z��#â�V�pd�gk�����N��� gV��v�bs'�o�dd�*cO�It=�.�.��	�L��Ǜ�Q>����,�@~�1�ItO{φ��wĠ���9�b����6�ə��J�_��N�i�\�냁
�,e[Z�����0�_(�:c����F�E���t�i$Ք���Nf�P�9Hc�b@��=o���t���
�����푹l�A|oS��V���=����ثm%a��I����-H�4:Hi�_!���Փ1&���ܟ.}�����y/W��F��ʏ���������M�Ĥ����D�%}�S��TS.2�+b{|�!{�%}������	�
9��x]36P,�G`�D�#��N�t�m��5�Q��]5����QM&W�@o�Z2At��qn(�@2����%�f��f��(�W��/aM�����ǘ��15��ux06������˙�Z΢}Ϗ�,�<4�JE�Ӗ֜4^���b��6�2'�d�f`G��Z`G�|�L�5S�ӫʏ�_�M_��R���`O���9�h�O�5�R�s\NV&PkW�kS���N�\]?:2?�+/\\���r���*���*@�#١�򳱳���ԸD��Xr���8ٚ�ǮH3��0�)�-*/�J̞]b���~��<�i��(.l�r�͟�d���Ł��w�i�髶`j�f��*��<ZJ2P�<�RVX.�U2���h��u)7���to@7�{�^7�%~�`�	@�51��t[�?qr`�u,y�%��N����ۣI�g"�����6�~��d��HZcoY���.�S�t�k��8c[u��ڀ���r#g`ɷ㥙�~[�0v�7)��� �d#�ҕ$�q��C���h�B����+�(��o�h�y���B)VXj\����9�w"O���b����Wy�RҬ ��\+^j���dhb`4�M?��I��L5�HE������쏁�m1��ƴ���ʄŘ'"T~}�}�8��IC��z>׊�dk�d��|> �g�v]�{�>^F� ���S�_10>��]2����W[�Kz�U��U��F�l�J��)��I��3����+�'�����Z���̌�I�J���R��+h��ѓtR��fR����}z�)��,Qx���@���G�7Ya�}�N6W�Y��䟢�iq�
��gBw���b��C2i[�W6o�����@~� ��Q�"G�k�Kl1�m���(e���
L���_5��.���&,��7�ud8诼dE&5L�`@n��]����ט/gI%9������k����:�f�˧�a	~��(.�����us��t�(��O�:C݋9�~�1��8�oN��c��1n����� ����ʚ�]����"�z����Z=/��a�ήYq�C)����&r�T2�֟7�O�i���[��Ն.�څ�1��zV�k�RR���q���!mN�l���Ƶ���*�4�s@1��̬�!��E�z
���@�N�@V������*1�]��Ns�N���@�X�tĞns���G��@���~9r��{���Q��Ú�k����)�N��M8U��w�h4������$
;����rM�쁭rE�#p/�\2I�NL�� �7�K�^_@t�}dpދ�a��� ƒ3��1���8i��%c��eFơ�ڪ�?b4G;d�b��"�sΖF�������~_�X��X+���E��_���î2*��%���)ub�#%\L-���	�e�jK"�$��g	�����t*j�8%�i�uq�w
�F�(`r�Z�7�k�3�����c��������YF�⬬���0��z�%��pv����%o,g�>�.E���;�"i� ��֐�9l�n#�����o��b4R�؝:f�[���B6�5wD����&!!O�
D��U�s$�Gg�:%O]�M���ΔR�ъ���*�[PEc�S芃���r��)i�|��o-Xy׸�8kf�C&[Tf��{����}��Z�Rg7�n��i���l\(g���Y�=A�hD���NR�-��J]��+oc���V�zf��D��$2�X5�����<�X[�6�����=ib��B����$j2����[a�i�N(fIӿ�f��}�L����Bs��J�O�F�SwaW5E�,�������������v��D�L{�P,l~{�{���}rP��e��������	��ZX�B�F��;���T��]����Y���	��!����Jo�>؅D_�>��Q��pO�`���kKV�ըl�QAcҒ��N	�*�H�?J���o�2UbX��a�F�p�`p��	��4'gB(���4��p�^,�h��Q���~�����+*M8+��>!ƭ\�$����+V�'3����ѦGCw���k8��ԟ]�|Ptro~�cѰ����"3QO��&�h���F�i��t_޿Y9�N�γWX��U��n�xJ\i������������&)ț�Kr��u�~��/a{�-xSg�cY�f��������ϨU�aUϡ�d�9� ���i�Ǥ��g:b��rJ,i!��J5t���ճ�t�Bo��YFaa�����`��f� �	�� �a� �Jn�z˔J������zg�9�cjN��!.�z�-Q�s��f.2:T��
�xjH� l0��1�;~bϓG:��Ԑ��?���` �ڒ�|��N-����'��\^	���pI�+u���9�$|����:�mq��"�|H-2c�"�K��Y��+"�GgF��)_��˒Y���̊�E:�����o�#�����J��w��R�'8	eб��Ҙhs��V�� $���RNG��;� ��OZ�?g��<���$���xwH��/,O��r�D���O�Zc����FQ(����63z�7�e���o��6I�%.�@!7�v�3y���a6�ݔ��B򀧉h]ݬ~´����M6�4����&�����Ai�Fm97/ cd��~�x�8�\�|�)��E:��	&�~��Áހ�����V��$'(�[���o�փ����*|��)�\*2�~~LP���9F&A��=����Z.y����=�d/�-:�ʺڇw�kj3�$CA@g�>����ť N��}B��ё���?�8c��H�X�� i��vg]��Ρ�J�w42�xD��bmKH�d��ϻ�M�R��u��b�&�šC�g�{�s�<$,Q��l�;�J3��`l汚A%��z��=��`�Z���_����"���F}�����P(0v>�"g0��OJ$��� �����o�\��ŦB�G��m����r�Ie��v�c!�!�}_�O^�2)e��~=�4�P���Ü	nR6�X��b���ߎ��U�WI_IS�	����q{ֻ�2��<�0z
ŏM[E�21X�3� �*�����8P�b�4�}@t��އ�p���)�+L�߬��ɲ���ԉ�]e����=}������NTg�%��=�X�_M6���7��܊�wq��i��M�d�����^zM�kKp�a���4���Ř�g����}�s�o�"޲U�"q�	�Ɩ�;@]L�9H׊7�2��i��;E��m �*u�N�D�K!w0*@y{�|���D,(>r��ZHp�Eœ�Bw3�mi�wR��CG�X�#��&��hw�J��,���)zB�o�1t5�6!�,A�,nU��� ��a��6m�[2�`N�ΙU�ؾKJZ w�R�gAa�V�m��U
���ū.);A눻��OV��j��H�A?�ٟ��*Oձ�yKd�F��3R��E�{�'�z��l������rea)���.?<�QP�O�XpȭnS�g��')Y��CpL �od�sf�O�T0p*�Q��p�"v���P�*��筨��,��Y�iA�7�r��^?���N���@7�3���tiv�$
�ɂ�M����8�����ʱ�Bo���M���4z���ӳ���h�P�N���"ܯsK�q�8��x�Tf�"�@�*"`��xܳ�w��cIV<����S��WW���?!���vNrYTц5�(����$]��a�`�{���6�Q�����͜��!��̠��Qdw<��b�q�/u���Tt.��u�q�y�m����u���žVȵ��[AG�1ZF8+��C�ِ��]��x�Ua��qLtթ��:�~� D��^����D~"���sb����Q7v�Ǐ���O��b�����R	�;^cLA����:�Moj�h	�j��Q�
�u����1��v����f��׸߱S��D3��:���'�0�o��A�1�bJ=KeC�W��	��Ĵ���y�'z9��/_�	�	�?�?�"vB̙��i,�Ci@���b�H����?�A�R� ���H���%��e����|�1e���9-*	s�,�k1�$�7$��T�:��sI1h��lbK����C����J.D�l�6��ϒo��_����`z��Sdjr<��nzQ���c܂��>"�>�:�b �i��Vi������M����T�P��-)��!�v�n��e$��M�<���i*}0��Ćߞ�͠n���������E� � �S�j��ŕZ��V�a���Q��4�H��/�<��W?���d�j!3o�� ՗�d�9�Q���h1�l�,㐟�����K�u���uG�D�iq#�q�|��9Z�p7���'HC?uE||.+�9��T�	<r�Hu��*�p�T_��B,�a?L��wUe{ٜm!��,:�0���;���>����q��E�>H:&��s�Dt�n�uY�B< �Ή�L*����dZ�S���[ΑT��MWw��Np.|����]�eż��}٢](|�و�������b��wڞ��GK�QSJvwk���j��S��F�S#���<��w��Ϟ��>��J�$A�[���o-&Et'1�J�9��mQ�������ɩ�6��D �Q��+�ѡ6���Q�*�1J��������Ȝa��X�jD<�Q�uWUu��;������xk��a�~	���(�/J*?;���A�@Od��,m,/����;��4��$���m.�q�^��.�Dn�B�QRh&zi�Qo	��q�Ɔ/(JK{YaA#�`�sX�ܨ_���5,H�-�����ER���'i��D�o����­|�(@ɧ����%a��x�=������W˷�f�$P����4j��2�����l����~+���Z\W���zQ�3�>�a�E��6��x#�kg�{�#�j�,\�%���@������|V;2E�60�r����B�	9���[�ں��,a*�)�^�l>���^
�l <��P���z��I�	~�/�EW��/^�U���A������f���	�x� ��oF{�gi�n}�x_�_ǔ�@��G�Wka26l�Ӛ܌��v��TI���Lqͦ�#:a��`�SYR������7:��3_wu~T�
��­Gքk��OK�]\ۯ��A��5�ګ��6x\����(|���pǻ�1M��ix1(SΧ�ͣ��pCBТ��	�G˙TW;�] ��;��lH�0�q����x�`|E�ڬT��'�t����w�ЎXq ��|7x���S䄐���e-nn�<���M�xxa��Fc��X��7ݙ��c�ͽ�{�@l�
rsoWW�&p�D���?�̾N)fw��b9�﮿��~�䍪�b�ix���{9�`cN�B��ʘ�R�)/\���|��0)A}�ɤ�@�q�D�.>�M2)~�4\ ||�/�����HD"�7�˚m� ��EX�[:`t��^	K�].��M��!Y�޽ӛ�h�\.�"֩t�9�]�"��Q�����j��|���I�̢3<�hQ Ꮔb������
�JR.�i�}���8
��\�> H�RV��F+��jر��I��uϺĐ�u��/��Ĭ�[�W���F4ˆ����:�Q�2\��@�)���!^<��"RL��Ы���܇���;�;KDI�X�+З)=�f>@�hC��ظX�[�����h��Z1��5Pqe��坛6�,��@�?
?����?�&��ſu���W��������1�w)OV,��p� "M��E 3GT�7{��[n����].�a|P%.���$	OL�&V: �|_+J�M@��k����(�ᕦ<���[d*0, +3����}pK�%Z���X�s����8i��+M�h[�D�2��+��@�@�pӀ��h�	'�ٜG�l$�)�(wo����#	G�0��'u*�@Q���9�<Q� ���}2F�nT���Q	O~s���P&?.����E��=Ze�|�2i����#5�oe�a7
����l�H&�mS�a�?�b_\g�J+L��Ĩ�}�r�7if����P.�b_G�2��_Bґ̠��mlx P����!���~l�e@l��O���͝M�O�H������b�F��ּ��m�M�G�艏>�a���`�O��-]��F�QC�4� �t%t ��`��kck���`�O�Ұ�����ܪ���pp�wo��f9�FE��C2![�鞹�e�����\<�4݇�hl����};�~�j��[�����o�tTl��E�Yݽʭ.?>o,��vn��y��i�8���r��&�*���F���՘'<�=�%��i�w�@S���>� ��}<��ޚ!�uZ�M�})Do%�+� ����|S7�Y�6;!��<-Ԅr��t�kȢ(�h��ϔu�v�Ӥc6�\_��j�+���po^[����]9R�ZZĹ��e���N�?�L��8�0��㵌�H�Z���7��d�ɻ��_�R��)t��+\���2h���(�xL�dMc�B3	I�j��X�uQ�ܠ�Қ� 4��0�UB�2�/��$1��k��E�V�(2��� �����4�)ʜ8;�,��㬉��L߭��Z��]��
َ��2��O���e�����_4f�TbU#�����~)�	hJN3ō��'*����/l��d	�7�����I�a�Y���^�sAL��ݏ�����m�ޖ'Xs����֡nI�\R�[�|�V��Y�j�1��tT�^<�&tI�ޗ>gr��	�ӕ�'sU�.\j�g�S�]�=T��T�l�o�� (3K+�&g��&�j�&	���c/���*nX�y/����}De�l� �j	.�3`:�{[�q�P�?��4IәRF]�i�5�f!L���e��p"����!vf�zԄ���>!��&��@=*O'#��t��z��h��o.S�q8Z~y,��ݧP�����$�Q�4gRq�4���+A���k�6f��F�VtR������&���d㲁�Ć5j�^ke��{��ت�/k27;�s���)u8$�,���������~����'y���9 s�l�.�p�@�Ϩ<Uϱ�}�3s/׏�h��+\[�=03�U��y��{���gb���5j�
aj�F\��ɼ�|T����d��'dO��UP��e�{�=�F��*����n��D�3���Tl�Y��1�^�	d l��m��]`�+O��x��}S�`���Fg�j���~q%{�����d�>)�(t�kԪ�����s>ê�����#�S6��~�b�&��<��uf��\K��H��`m���%�QY��)&��F�U2o�zi�!1�T*Bj� 0i>ڮ�F^��(T�
��T�ո�	�j�.ǤU��W�׍w���/��c������R�@��b�{����le�w��oY�Q1�3W�'.K52O�:�i(�u��`~:��t�����
�R\��N��'�J�"=��[�f��TG,�g`{����k���%3��,��p8�L;��w��!��~�@o<Q-��P��={�h���R��'�FҖȸ��%Ŷ�`cf��*&��0i�U���渁�'�ˊ�,V͟�!��=M��GX�<~��]�.m}�>���Z�"��<��\�f�z�������
D<96�,�� h�V��:'z�9*f梌~ޡ��z+)�d!XW�� ;4n�G�V��� ���5�ͅ0����ᰜ�褊˫�ll�6�i�q�	�w� %�}z�g��sU�Ľq���>�.h�Q:������"4�U�������!P�u7���w<b#Q�������5 ����ؿsyz=�#����W�OWY^U(�b͔��	�l�b�3����E̹x�	'ݟ�b�]�O����\��vBx�hX��tP�\\9:7�m��r�al*�*j�9�ᡓK��=����<�o^)ݷ�m�������Ѿ:���a�s����f'�SqzH8�ӈ���X9v�Dz�Cv3*�H��x���b�^�I���z`ƪ�i�m�6�lYo�5��|�v�u2����{�\7�m���Kؘsa�t��yC1��h�V ´�HQ��#i%c����m0�<ǭ�9�"肕+Q��T�G%��S�Lx-HNw���Pˋ�<�J�������%t|�P�R@�Gk�,�Azt:���}�����
J��|�@�"�Yq�W^@�u�z����Y�=/v���wb/,���R@)X��p%�(U��"G#���[}�!-h9��WX3�:ŭ"�n����D+�#����}$M���|���j�#ιI9�R��Н�fm�±�|��C���pPdWN+��,rbs�VP��q�cx�uY�k�ƃ�_Y;#q(ۗ�bh�t<6[�a�G�!�C��5�cI�ɒJ�U/dY��{��e�&(K����r{�7'�=���Q�P2����z綩.�#��g��n��o5ʒp�Zc�����	b�`f3�TqT�ټu�Be�%tpL�0)������:JS
�J�?<~O�C�dt/q�\���ܝ�ˁh���a]��d��Sc�,�j�=��ikM��*��#��f�g����`T1�e2���^���SH4D��XW׀�=d{qN��{���`!����'+Y3)~�}p�W���[2��Qnv�Ig�e��9�#5�Z�+�������@�Vd�y��:�"��i���v3���ٟ,� �S�����n�&�t(�v�]��<h�^��vE���a�X�I3�v�.��Z'^\��ާ�b|#���⺄�����FqQʝ9�!�Tԫ>D����o���dj+�f�p��������*��Wo�|$#�(�v��&���{�!{�r�,�ճ�5k���C���ށ��&�z�o���X���;�Ѯt���uc���w�u�9�a��i����6z�+AԌ~�^�Z�\��6S�lkHw^{�>?�g}��=��oC�R��Bc�*Ķ�2ޖ�����?M�0d���R!�F��Uy�TB��I����N!��]�s��ej�p�M{w}�낫�� �lf�D���u�ѡou��v�/� �PK��p��	��0�Ɵ��a�Q-�ޛ����>n+�+�_ZG�f��.d�a�~ba6v�0l��TN���cq��$�*"�aGp�,t�������\���k�sdX¿�b��;%X��_c�yI�uLm��Bp#Wj�6]aon�f?k묩�Q�z�����wM�2��QjU������ȓ���o�ѹJ����Ɓ�>:��v���G/��#@j�\#��*�T�2�w��?HU�#���"+pk�CӖM�rC<�͵��`���5Q�5�䰫\e���(�3ԗXÂD�"֮4�ϙɬ�X�mAy=.�z�BH���EEd����h�ػ�qY��|#����%�\R��QG��WN���3{;,����ix��@%�)�N_+�Pn�T]j�e����<���
���#�JG����f�C�c(�װ�!qk�\6��'�S�$A)jSV%�6�/�k3��������G�n��݊��L0pHC��R0�����<
SB���iqۃ�_�>�����k�t1��I�q��]9Pv�����K#��UϽ

V��ru|7��EI��ژ"���D]ʟ�9��B�5b��n�C^�S	)zu7ZX���p��6��$'������)�h��Zr_h�[EJ����dD*�9��ۮ�TLXw�D��ᰲc��cO��H엔gF���:�lͥӱې��bb���ӌ�ۋ�9n+�3�8��B]���[�Yy���TQo%����F�^�҅>�lFN�q�����[��(�z�2���T���w�cr���e�����w6^z�w��`��]рJ��P�F�|�	�^��@��Y;�CS�<<t��#�x�������艭����z�`���^�W�}���f�-�
���+/�N��t�w�"�(��5�D|6��ۇu/ױI��/�u�N0X�_�O��fƕ�Ou�8z�������2
�=Y8eX�~)�5�ߣ�t�<�~K�Lqv����D����"D�+�aMbt�"�ѷ��%��"���=0�}�4o�
N�<�y��	ksf��S�goO��=��J�P�h��DL\2T�����xzO�������Ԗh]�U�Ǽ���Sy0��F�Ic\U&������iL����tm�f�[� 秡*�D�O#�Z�m���Ǡ2���������4r	f��p�
n�Ǒ�[/���S�S�v���ݚ�(2�X� ?^���ޗF��թzv�i��`��0s�:��t��ĝ%�:���R-�z�J��F�'�6'�:���z�~�R�_*/(���:�+Qï��������rX�,֜]��90����6��<�w�o��.k.3p�׷"$��鋒�; ����r?���8����u�����,���x���or�;�*��м!(#��{��ނ�:���.�ׯWH�c��.��%��'x-[@&̪N�8��.Z*7#/��Ee,�
g���)i�t�F	�h�8~�RLҁD��yRq��F1�q�#3u��f�g(Fm�$9��b3k��H���T���].��k̍R��//�a�6)��#�Q�'�r}Oq	��3`�rԤzŚ9��V<��?�/}�0��E��4;F���b�V�l�VCc��`w��x�)zVx�l铭����j��6��6nsń"࠭��nz9*z��N�w��\P��Ip �q_c���h|�J��i�k�<=6};���i57O����(�pr�ʜ$�b
aRD���16�����!��rВ�gB�A_u�|��_wPu����#�e�;���d�����B3t�X�$w�\��vVCǂ=ΎB�����F��W��>�kU6�v�O��si�4{�s�d��4�%��q��y��&Va���i%�m����ï8zI��$(��ڒ3q�3���jB�2$��}S<2���.��a�,�l]��z�6م� 滩��A�';�ժ�it���\p�����5�w��௸>���6Y�{3ᴐ����դg�u�#r��7�M!��X���㴫�`��|mX3���z�+ٰx�3�jq�F.��i�pPb�cbR?�"�{'� s�����s�Gi�'C�����,�+, �XF�e�����*y" )S�,҅����񛌂��������R�9B+�c������V�������z��=V��k��%��l�5;�mU��X��I�9������C�4�F��nZoٝ�6u d��^��Mf���7Q%�k2eu�wP�g���%�2&I��gwǹġ���*�v4�/���N߉����2�d�l6�Y��	 ���-�BI��4����q_��"AMY�]�s�:2�����V��LOgt˃���J�����-[��w+oْ��U ��M'��m�>�3#�?�0�FPXټ6x |!	ֳ�m�2H�����h�b)������:��Z���v��`ԕ_{��2߰�|� c��ۊ�ll�}�!_L��j�h�' @G�/k:�1Ɨk������!m�G���1�		�t}5\�����@,-�^ß��/�B!V��}��F�����X�2��73=�q�0��v#��U���N�k8<��c����v�KZ��,r���!�W�Yte,��5�â)��gM�u�a#U.��j|@�~���׺�a�x
�*�n�?�P����V��lV�u&�Q�?Y)�]�%�5.5�,-����ذ�}O*{|����-v�uG��,o�ď�q�~Y�(U� ��c#A�������}�ꡦ.?�=�篯Ta� ^b��-��@�R|��}��b����p����2�#��! �4����+-��N�]��,Oa-G����F��0-x*��N-�MRR�e<��*/�\}J.�vdi���^�]N���%�D%b�酝�g?s�@k+m��K��w$M��k"�lP4n�O	#CV���i�Ùu���������F����v��y�c{��25]��z����,˹���DD�{ѣ?���x��%K��Bnz�hd�/N�����!��"�L4(8�<�p����h��x]/����������m�\N�X9�م��^�Pq�ۛ�I(���;�Z������g�M��hc�����t�Sr�<�t�X�M�.����z���	{��0FqM�c{���C*Ի���1r'��¸�Dv��U��KL���v���?��7q40u�l~P�e͑ʂ��	�o�����e~�I,R���_c;Q�Vig�`�4e�V
��1Ċ.[��t�5a�������,Y*�
Sv�Cҝ�3b7:���s:�������[���e^�n�H.7�M^ ���n
���r�@����Bd�c��U�887���i��{�I���P>��-�¥7[TR i��3)�6sY>�y�㘰-�H��Z������F���}��PPvW�������%��6xֳ ]�.������U2�o�I��A2��KX����a�Ђ0�������o>I�@��}�7{��q�ݺe��o&��.f�kia��;0���[�6-��/��Z�0�H���'�n�Tu��+Qώlh�.�?�13�(���e�J���Ef돴X���C	�om���K�4��vkT�Z��HUk���;|����f���[������uT�0�1^��[�␘]��s��h�-<j���G��S�?��Hlb7����7kޅ�i�ܘ�+���v�{2��E�z�-��U⊁l����#��d�r�;"����"��{���~֘�Q�{󏼫�'�i����* B�B�;I�P]�8��P��
�9��:E�Vu$|Ґӡ�{<��_�V���5�9gL����3pM_�L�id?�<1�;5@@a5���2�P��Q9����_*�E�����T��~74�Ν��$�i`I'�;�r��@j�#W��.�%����{2JnK�zN�s�����O����1�i(���|a����K�D��J�Qk�%�\ORN4įQ&��Wv�b�P�����Ӵ�d�E~�[�����*��@w��_���_ig�x3����T#J���=�..7� 6�����N�
��M��H ��jg[յ#�`��?��M�Be;3+`�q��l��S��8���$U�ﴽ�z/��F�iN�~���~"�y��)�w��X5�z4;��������fT� �̥����m좭��26�.��'�Yj<�N��p.HA�Xg��u.j�`��~β7�3��?�q����gӨ���l���%�w�z&��l~pz� h����;��H�$؎L2���q��XX�s9�+x��n*�?v�ss6�v(i*)ϯ��ʷ:�>�^;���%� 5ɡ0��08>d%'��T�S=�}}��<̵����"_J{�����^KG=�Pl��fɲ9����d�(�s!���l����S��q�T�OAy�����W`�|?Xȩ�������q�y�_�e�Xr^�ߚ�'�nL��R�g��}��m�Z�����.��ʽa�SC��H�q�\ �b�ty�$'z�i���#|�6�81�Z�Ģ��.k�.ч�?�X�rxS��}�]�T�2��bo*9��?u�( ���V}�o��q�QJ��?��|6Ca��P�!��i�QC|��R��5�̻�&�SF�XAԉćk𓬌�$������#��Nݗ��`Ĕ�u���i�8�kҵ'a���o�cb�@ްj��I�j��"�(�h�\�ϛ�v����o�&M�� \p���kVz�_����V�|x��Q��׳n��_�)��$׃��=�k&E;G'��AMr�~Ci�Ւ��5��W���$��H��{"�(�Q�g��Xf��QcE2��τ^/;�ш7u��f���ɋ`�z�ʡ�?�Ծݵ	u�$s��0���8C�9@&��:�";(�/P^�V�B�&�h�����$<
�R)�F���`�7V�DOC���y<��ު��H��P�Zoq�ׁ[�`~7���*���ک��R�J� �r�Xg�Oo�!`����A�?c;����Ddrp3��J�@4�&F-��n��;�V$���/�Y-/x# /�i�����䜧&?�hX�]u��ӣ��Y`1���XJߊ��"m�{H���yF����SQ6᫫(�v��	�/�-�'�g�)>n�Yw+[���I̑�A��ʖjw<mK/L{��$�NԀ��uz)�t��>�Hۤ�>
#��7���G��7����2-�R數�$���g�*>��f�"cR��sҩ�4�5���@��Q�}P�����ϲDU�D��U����^��Znʧ$`m�E�fN��P\H�x��A�c��\�1ސ:a��`eC���]�֘���ꥁ
���e#q�l;$)L�����n�N�Y�.�����@��a�4F�ojh!�9�h�Ǳ��޲�����l[�����6�F�ϣ|���%V?.`ݞv\�'��e�?z{�[gl�u��%K�1�Ѳ���H��uu4+5[.�m\��7�g�d=���I��p�PKso	���Uc%"��kiQ��6�vh:U�l�K5mW73�����I��;7�.2���(��P�&����>�yO>M>�)�Z��G6G�u�����Wz�X�0�D�(��>-̍{a	p��G���a)�����?����mH���aa�5�9/N�4GД�-<J<Kf
v|�'Q��0��4��D�'6�f]2R��;�0o�
�E~�>X�WP�:��_��7��{H֔	FƜ4�O��YK�\J6S�{縈��a����� �?wE|�@Y�.CX�ze#k�<�y�S$��L���B��,�V��r���ԜH)�C_���S~$�E��]+z�=��[����**~�7����u�U�U���o�P%ea�����D-& �gO v��+y'����^���n��*gǋ)��>��E������ngB�E�o��X�{B��a��h8^A[�+45�\jl���ٞ�cB��/�6[Q�ϼ[%��dN�a���,�J�ڨâ�	;݀;N��J\ӏ�?��s0�t�z'%.z����<�`U�:��1Q�z<]_��n��lٓyP���>
c�tRy�Z�h��{f�n�������E����֏?��;D��5&a�t�����\�R�,*�-��2J+�^��?&�2'4.n!zw=a1g˕|�a��]��{�o�iow��k����G�W�;��0�8�k,jP��uN��lO慔�G+�����þ�iw��}����	�V�U����%o�[�����.����&WP`YCo�$�	�\����歉&:o&$��!g�]C_�P�ֺ����u*C�b�a�rJ4�~qX'���|A;��>E�f<A��i�r�dp����_bF�:v6m��ё����#Ч6��k�������|�5@�����}����C�z��O����f;��������«�(���������[�h��k&F�@��?ͫR�lC5D�~'��A"4('�ń���0S΅�o����˷L�����k��>�waS�N��L�zp� ���z�s�6�s���a��S�4P@�8\�8 ��5:�Z��'�Eo�/	�K�γ�[wJa�����&!���|�g�.	���LU�	t͝�6|}mC�j�m�wƠE}7�����6$:Ư�!LN
�AU���~�G���8��[ꝟ�Z���fw�b�-sp��I"� !\v V�j%Y�ך�@�9���!I�h���8h�,����M��F���-���J����N!j�/��#��V@r?۝�T(�� S>1ξuA���z�Iڳm2�ֳ"J�#��/z��P�M�E�H}-h�9�
|�J�@�xH<߸�(��I?Gy����bӼ�ejGe�N�����h�6l�c���
�V��K#}���dC�n�8
�\k�e�c��n�vf]t�Wu˃�(�ɥ9K%�ۺ�_a�F��QGԩ	���݉��n�H!u�r�e%:16<�қ律�e4�+7o��7�WGJ�E������u��M�˃��tV�PEU�(��u6�hRÕ���b'Yg���i݂� 	;�د��R=�c
��or~�e��@�N��Q�ݎ�?��	�/��&}c5S�g�[U{*8�q�[�G�}ӕy�7���`W��O@\�XVיpHs���n�[ �.)kP߈�g �Uḅ��Zo��~@+l}H bS%��M6���R1��!�O��p��1���w����w8j��iD�*-�m��ٟ0n������;^J~n��h�P.	t��]� '���KT�_�g��$?�S��R'��?j�OF�Zt�@o�@�aQv�����*���[���x|	�t3��$�c�6͠����Bp0��ɋ!`��}I�$���j+��e��v�t�D8�#�E�AH���:_̧�Y�Z�䲸=���9έ<��T��lxߎ/�f���yt����K�넺���E�%S�1O���Q/�B#K��/�^f��87�3@�iti0��;��T{��u0�ś|/�_�ȧ�(�����@伀�'���@J��G�$�"|S_O(�,i���bo���ɧՙڈ��79�&[��{�\Wv�����~�>��-8�����d��|���xZ��Mp��n��k��	k�'�pu��W�G7������:b�:��%���Q�c����ھ�nò���F�r9�Od����,�NL�>�����_
��}{7�dj��S���(���W*�u��9��V��	��[ҭ��.蝌����L�����0�B�h'��K/&��8��b�Z
;�v4(��d�s�t"�a�$�.p��R������?��3?R��[]�QU��
����F���	�2b�C8[���~Y��Sml"`�3��;�W9��.^�Rs,[`H[�f(���y�$���¡#M�-�R%��+�n���ݹ�f�Z�dssRc�(wn�@��у�]\�c�x�_�S�_.�Ӭ��)j�y�Ӷ}��N H��\�cq ��e`�VeDx�i��bX��W�R?ݱR����{�{��n�*1g��7�>�k��}BD��F/8M��bE٨yˤ�«O�'�a5V���8nC�V�1�����ˤ����~����m�a�S�3���pF�:$]��Cj��Pҥ�W�LX��N�;9$8��d]��v��>��lNWJ�#u #@U�EO�� �7X6_&2߶��%i����M�a�s����Q����xJ	`�T�5��rچ֜EL��mk�Ʈ����.R�iR�6���j�o&�S���U=�
IUOb��d`�J��{8�K���{$��h:�}@r>�1�s]L͙� �m��|t��i�����uM����k��֢���HE@+��~Ɲ{�z����%��D���|�(h��Ǌ���.������:����e�>���+�~98�ljjz�bw���?�Y@���� ��%Zh�l�.8 ;�>�B��>x3�\2��+� ���5�8n|ltFP�։��&�#�O����]����D`$�Y$\3fL}G���az�l��U��z*��-�~YE���P�CJ~Ř]r�0�Y;;�C=2������+�M�F�++�sE�S�����,+��s�����i2]B��M�����بjM�ր?*�:FF�>�;��9%�����;W70���'7}�)��A�F.�^��Ҫ���r#Q>9��\�W��T.���L��u�R�)2,O���B�ͭ��ָ��A��=�S�.S�/���
P�`;�zI���3]Ҵ��c��~���%��W���������',p���R��qEQӕ����iO?�h:wϵ�c����1s{}��	�_`�^D�U�]��J8f���e�fF��Yb��9U-��j����d��1���ἇfr�	�2�Wh�w�+���H��\�������	B�����$A�F��E>8�/���.��&�222]��������$n=�͒��T�A �R�/d�X�f��M���`t��+g�0��T���!�sDc�ld��dG՗Ӑ��,���fE$^UZ��T�6��k"��.�D1�7���0��d��˹��s��������4]�ݧ����$��H�?�X<��m�Ehįˌ]F�8D�����L�@�9@��٫ZI))���4����F��G�Z��&�:��oNsE%j/�1
��� X���p��-bx���z���k����g��q�"y&��݌��Ġ���μ��PGGˡ!M[-P�m1��`r$M�=�g@�qj=cӼ�>s�b��Gx^�(�<m��E�B\�Y@;�[
h���fO̹�w篱U�y������9`�����r��yb>���6�;C��G�%��	���j�'Qg�WmS�D�kӑ��4��^�R���0JO�zJ����H�텙1K����w{��I�f9q41��|���+��h�gPD���92�l��m�W(,_�4���]�ޥs4�C�>	�QH*��:��9�ɑ�ւB������U�v��Иo��#[h�p���I�2;�Ȫ
�3�N�ò��B�y��n�9�g�=3$B$z���k�Ԟ��R�K�tH��IO��)|�=\���tE�cu�x�?��v�i&.�k���*�gm���!
2���AX|L���3*�сțH�gm���� �R�T;c���`�
�_tR(�%������f8����,�~G#��">lß40��ʴ��˕0;x�1%�M@�z⮏+g�U*�4Ғe=�ÇL��kjѮ�$�蘦��k��	X�*F��ڒ5H�x7m��Tr�tϧ=c�fXߑ!)�L�V�R2*<��|$�G�����1K�>.���ؕ��6�ۂ徊��qx����CC��Ե$�9;o	bV��@�Ti׮���g��j�b�g�f؎,����3/�<��sDw_��f6"�)�yPri�� @�2`������CD�!���|���w��A`*�b��mTOs�/�Z�v�=��ME{��&����ng~�)Π ݵ�uՒ�c�t��T	p�+h�&� �H�ɾv��_x����1�+�P����T��>��^x0��m�����Vw�[�Ġ0~�k�6���z�?�dX@������F�7�:΅ ����ʡ��:R����)��o#Gt]�=�~?�;�n� "�CA/�E����"���8�G��*�%MAü?���,H>dؿ����@����4�� ?�V��")��n���&7�Q��qW�r�k`�XC������k�m�@7-{a��l��JJ��p�I[mI?�4�|�J�d��y�UI� �|�l44�H�8Sx����C���VA���NV��?R�G`��N%���=X�����Dl\���ɿv�	��n!�6xd�Ӫl9���C��"b�;G��"o��v$~�:n@�>}�2��L��nT�u�&�8��M�Py,H�x���I?��VBc*v�V�in���>{G�s�/�)(��
���?+'iNｌ���\�F�8�5�1Ş��e�JO�{���y��2T��<�Ɉ�G��@e�`�u��agrQ�R6D��&a�B�A��oߔ�!�'�V����;�{,G��{pͳ�?���ʞ���Y���n��-�B�����:��G�^�����{�q�E����B��W�G�F��o�?��	+�L��v8�l)qh1]�Y��Sz5Z�>�u��Q�乖y�
�$����g/�!+�i�;�kU83ΌL��(\H��2�k`�-�%RWf�Bh Hˇ#�ן�! m�?����R�ͫ?���Þ��{<���N^�z���!+0dM�%N��=��;I�x�t�s �2@�Q��K�H����a��_�Ѧ�kXa� �ِ]H
n���紦h��e[6�a3�0�.gv�D�Ҭ\��#�̇�!�,^����Gl��~�/9a���r�j-5�hTpldZ�����gI����Y�=���������1L��K>�=�oKl8�S�Î�7T���@�
#� �C���&C���CL&-�����B��*8�<���5z��Wʊ?ρ�'(4]�p�3��-A��\�Bb�z�?�D�w�~~�.��_�	K�Z���Re@�|�k+�KS��O�m�Z�ԝ�=f��(3�Dv�1�����iz�]:���X����:��p�
���Р$�:w67���㻹"�E$�)Ԙ��3?���}��DZDE+aY7}��;0�dW
�#g?�q~�����,�=9�L��/.��U�\�=?�͚î+�}dU8��9�	W��-_R��F0n,�yuL<ND��O���Tј��=����8�m`��	60�kӵ(�т�%=���&�I���W���n(Fo��w�y �G���oRvlI��Mc+���*��/�F/����GF��J�e�B-m�'�W��7eH�X]*g����#^�օ���tí��^4��o�1If԰� �K���L}<��  �?˸wAmj,"��1h|Bj=׏��F��}<I�n��^Z�>"{�8*����<{����Юzm D]q8F�J�r�R&L'I����H���<� 4��&�Nh��j�e\�����/��@����X�� \v�i��k���نϺFQn+2<ۼ\���\A�&��򯺯�~��l�3��s��{ϥ�(r�Az����2Swˢ㼾9(T��$JnJ�.�@����<�1�۟B!���GG*:�$��8��v��l=�E�~X9�?K�̜^{Ƚ8������+-N�~�*Ɯ��;�b�����T���_[Qy�;!fi�VH��{`#����[<�G]�9����G��tY����q�|ߓ��QH`D�e�,W�1m"��Q]�HUf7���}Dw���>�8)�����jP�?���Ξ[N�!/��0e�~�WƟ����_�є�Vߵ�'�ږ����Ʉ[�]x��ו���y������rS+;�;=uӇ�MZ�<���Rk�U�ݤ�%�H�DXf\�#�FOb��S��z��:zj/�Jkև^*������U�
�='�qHI{8�h�Y3(ܟ��,J�U�ej��L8�_��F���O��R2R�sG�g�җb�� �Y%�G�ň�\X�5۞�ǰ7�=�	���G���޷�4U_�a�p�ѥ�#���y{��rr��Z���3}2�z4������	������|��<�5�w�L�v)]��2	�͇[�cN�J�D���n�
ׇ�ѽ����S�͊ǣH�~)<j��虐�F)<:�i���i�������k�ԮX$�*��_��o\l��[]_9�M��7����`�Ax�������	��vҲ&����a�{{�Xqt��C���:0�W�Ά����6~0E`,��TZ�0��������<��(����i�`��S�����z{A4݁�T5��2Y��o��e����6|����A�:���Xu%%��Ӯ9 *���C;Q�
�
�y� u�Ͱ#e�WiЏa�9�g~�����zo�Z\�m��#�1���=��C�s����×n[B3Ǹq���h7��MjzY�Ai��؆����q���0�:ť` ��S�DH�.�l@����>���~�H���,yM�@��oE�����S�{�5],���8�{�zx�i�trE��|i+�|_�Ԭ���8oRz�����64��(W��6=!{��I5|�ݚ�� ����O���%5{k'1-��l�Uj�](��Ab(�0�@�c*��VM�a� [��kh�E3��È[��s��`���,��	��N��blTl87frS��;�ᄭ,/���!5)�!]��U8������ת��Q���6�25U����W����^\J�`~�_�@�&�7JQ�\��)�v��P�=>d�sc���}���/�<\�q}�y�+LQP%آ_mͯ�]TZ4*���1T�G[q�Ml��u�UGeC};Ta/�>I/���ٴ2����C�ߡ(ze:Ү`�Z%/�HV�
4(�V��C�r��;Ў<u�KbwX�r�;|<���n,�O�׾���HuN�.*Tf����AT��7��։>�IMWPC1������J�tmv�ְ�TYH`��B@�ظ����k%�wݜ���]��G�	t�imaw4�g����΢^:*��m���8�δ�ˮN0��J��י���ur{A�z�
Qyw�f�VK:YK@l= B�a�bt��*ú�o6�������3SI�Tܢ^��q	��W�󋅠����@�@��Z���k����>�r�j��@h�QSq�,b�aB ��*{�*��ϑc��5Ù�:=+���d�줍��+����<��㵵�����2���>Q��}S�N���4��FQ���^f
�M�+|�Zg<���eN�z�X`���Uw�F��O�K�!�}�"X_w-�_-1X\��R����?�"p���"�����{���> ��N3*�����6Lf6�lZ�<�$�y�[��#^ep?������/XY����E����2�|���_R�&���MיQ�A������_V�hN�nP�>�%�g9��e?�_Q^A������8�#��(��z�����G��\��̫!�s��r���.t}ɚ7���o�*D�~�k|�<��Զ��7��!9����'���
�D�$j����U�>:?3WA\�����<�[gR�����������	'��m��B�"3R̓{1u��EXY �;�����2��������>75�{V�FL9V���0��C���K���7ެ�VtL���o�d�	a�&x��V�5ǀ����?r��x�oۗ3y�'�N��I�p�e&�2��7a�\.~=w����ޮ6��J�􀑼gݷ�a�	�Z�U�7���m~�/��IC�eΗ(�Y����BA��S�����%+.�]�9�
O�
�w^���F
}�����J�lwg��>��m�ЊW�-�\�X<i�o�.�- ��q]*O��fɁ����֗�o-�f���#'d>U*�_�\_�����U)R�3侢D��Kp�IY=���/I]��p�b�P0�
 ӵ���l
�n�Ʀ;q�O�Y����vXX9����AE�zo��*^���}#�<�8}Mp-�٢h���
:�q{Q;��%�@Z�>ƥx��-$BY>����,6��O#F���`���Q!��[��aތ��Y�v��
!�i��4��O���J�f���w=����֠{��("���kZ��$��!�l�ZJgh�\���@.��>����(ɳL��͗�ܚ_�} � �RJfu'�h���?��@5 �H�p�:F���2��w��)��ɴ�A�]6y����m�.�*�1EԌp��
{����iDm�#Tj�T�f�/��6[lI9I�u	�t�;$1�Q�t���O�#�3���zZ�P{�-L�(U_��TeQ�1����P�}��حW�E��iޯ���k��8�Hr[J?
��R I6��?�2+a� ��wÿ�����}�f=!�;7�����I#�dZSQ�zh����$���G��ި�F˺�c(���m�BZ�q\���ษ���Oh
5,��`�A�����r\�0�`�k}���"03DN�3����y���GP"˥RgE$s@������"sT��V2�;�7��Wy{s���O�Iٷ��r�Ki�>����5�å.�S���d�犕�:��0{B�\�>�]��K��<�;���׈�i>���Ki\��3��"���d!�:���_�7�$�.�^�,i��:�~��9>�p©�RJ���������.�l�Gk�C��4
�Հo�aM�SL��e�9��H��V�K����Y5p���0�䩽�D5S������(�������Ϧ8�˽,�K�-#�Hڦ����[\@�%�W��,$��غ�sp�0��ϊ'���3���8ݱ�*	��8���]�}��sFQ�(�EqXzS�2^s����QKj�RTb5fdY��>9���$�C�'i(�ޘ)��
q��]X`�d�Ύd�<��� ڵb�x�{�5�;V�W��U��b����j<�B�f��|�I�h!q��[<	���Fﱋ�F����;;LMzװV���U8/&5,Uw�R���y��X��ƿKm=��{�I~����<����>�9�D
�5x�dCJ�ͧ���7�1��4�8�����F~����C{�q�Es!*Ē8E�T���ub�C�u�3��+qs�L2����i��U�qi{��Ò�0
7���	�����b�����&�k�T~܅0W���B_��H����ح�B�d5O�Yz�׍l6�W���)ϗX����2����_�!�\9��c������\�rTu��
���k�Q w�����FzN<�פ�bQ���!�ߓ֢�a����t�l�8��zU��K���HQI�-�O-��R���%���ϒk<�|���A��2t61^~�*ަ��2Q�{���l��H�nm�����}�9�h��+S;���=_&l9�Je��7�viRTNZ�h�dsaT_���b��������í+���ȓ����i���K�0��z�p�s�S�L�Do
	�Ò�:<A��\ڣ����-�\d��]�-t[n��!�̿��ݿc֝Mj��Js3]�X��i��e�����"+�N��'��kK䂷���H�{|�T(� �MU�b>VCڪc�5��.�}��y�3@��n�δ��>/�J�`I��5�x���# %��Z��Z��T���9Kc���D�{��"<� ʳsY�վ�_�8\���N�+��}o�� �cύj�1�ӈ<� 4�r7Ɖ@��:͸d`\A�"D]���0`{<��i���M��Aв1}�:.�"K��Ӕ����%|�-����|�6�q8��&���
oM�Tӿ�7�0l,�����b��4���\�B����ш;������t�X:�چx�'/\�]XA�7.� � #U���2K�grO��}`����p%Bɏ��옌�%PFW���۱=,tsB�(���cb�����W4_d�L�$���c�e�
�񈁀�L�xGа�D�u��X*L"�N"���6�a��!�c�x%Մ6{M�q��)�_W��ϝ����<�����6�B�ڽ��z�((P�m�L.��r��_F�D<�,�*�62�Q�ӆb�H�-�t7�/�;�H��X�j��ԺI�G��ܼ�ʜ[�TL8��y�K4�N��7����)��A�9N�2��(Y�$��u~غ�*$��^ě.�X����D�-�#��N�e���U�j��B�I`��� ��-�?��m�,BJn��d���:;t�!x�»�wX�q��Yo����J�h��9���[�B`}C��_aW�;$rha3�	�(z���cמNO3�� #crܽx~�9�$�t˳�����
&J���X�r:�O�n���v��{����<	��D(�n�گx�C���{���v�g�;��ij��Nw����Y���	ql�-a��SS���:��-��aS��~���&�J��&#��`��0�<��%1*��"W��P�.��*�_�+X�*80�,��YJlH�-��a1V;�$�,&E�G��������b��F̄�|�'�!����j�m�����Iz�h`����򞐕Aa0�[�V�HOLeZ�fI�'[#��E��a�s��s�Փ}��%xB�X���7e������8�*Ư[Ш����(�\���^����yb�ª�0(�4q�X+��:��'�sY�I��EE�3�,���������<��!������mP)H��>�=�̚<dW�_���Y>U�.�ZT��H"d�%H�r�_��wqr��Q�A�1_L�Oe�z"gV�TwO�'6��!�'�Q��T��e���8��m&F�Vv����N�=����&�"!�\Dz�-��'D�����u�:�~Ra�HP�.��VO���\�D�xbՓ@���-�bߕژr�ˈ�3G��|u�y�v��N�#>�Q���VT[�B�$�ƁΧ�`�����V%y9	����)�f�>̧�Ѳ�!.���;8%��ko��`e�RP��MmC�FI�_^
&xQo� υ��1�(��/��,��B����R5�_����2��Ô��ϔq������I�O]J��Ik��|������
H��k 
���G��3��7+qة�݋g�!$��-��F����*�"oא2��:���%��o4m�	5�'R�D֓�nkE4Í��xB��}�M���E�0p��I�t��м��������1���f����޶����D$u�m�Lh�����+m�p��� =.rӇ��A���F�q�3ޗL�H��=���T�P���`���p?�������:cUUʕl@(0d�G5�C��L�֘��.z2m��j���>Q�6W�A�����T`�C^�ofMRw�Z��kJS��y�_�P��{��ߠ�CR��,�62^�<�{*}�r��N��AB=݁��mVZvu�����t�&�(�MU3e���c��y�֪�ʚ�;
-�n?�v��`��hq�c/R�썏��k\�V渚��]�������#@��xD�_G瀘=M�\%Ꮚ3|�S�{�����=� +[ɼ�K��~��~���Qڥ�\7�ho�JP�P����NZKп��n�d$2�(e���д�0�]�ʾʩd��2��,���g!L'T!���tK̑`��ρ�t���U�DE�S�<[=������+�+�<��~�~	���}e�qB��oX���	��~�_M�ݨ�[��'�S�h��t� �_�KrǒB{��Ƹ�7΋ka�I+r>!���� r6��?\�t�ַ���a����Y�/yCd2���3��Q�EX�j6F"/V�a��Ҹ�tE�
k����W�:.�5�����s��}y�iФ�&�g{ �@����AVO!�2	���N�j��f1�����$Rf�M��Y�<�P�d��H�"���ܮ�	�M�b�)|�k���C��s�6�6n>�ega�9ĩiy�T:Δ��~�B�z1�y�������)����J=�L]X�>(��R��.��]��#'��T=�[�>Ezi,S��hO/�\\���\���2+Q߹g7?8�SS�i��N�j'$Y�)�gu���z�YK�9�0��!�����w���w��<c��z��r���|a�=Z\x�u�>27���9�E�����jAw�?@�����dT��]���N`C��>C[��O��7�*��R<�;HJc�Vgi�>�,L�<"�שnt���ءm����Ώ4�
>}������)pO^G�>؉��lZn����
*(C�ht���+b�HP>_9�j�*�̌sgx��l�N�E�'��O�e�3~�l&@xd���CB��gԋ<@�o �[�����6V��� 1[�QD�v�n��pd9
��#��$>�oW���,�%�+����� !R�'vxJұ�Z`R4ۀ^�Ġ��,P0�恠�>�HR�� �����z���v�@+Z,fpzf���8	�~�q���\j�L��f����}����/����Qp��볁)%�Mj��us9�uQZ;�!�>��#�2թ�ND����
�/$F�h�T|bY-���7� w�jc�a�����U m^���J��.����ʵԣ>�+MH�T�֪��� �-�OmС�`r4oP�&|	19�ЫoS �HG�^l��oJBT�&mR��j�(�m~�SI�_�Z�*TuN2z�o���Z�؍+��f�Lˏ��kfp{4)�M�����&ET���{�`�!���L\��N.Rh��Tz �<b?��ص�6���,�2�b�ĖY*�,4
!6��ޒ������⻣\�1�ܿ��k�񾏕�l���.!|xx�)�(�~|=x�0��G��"��㐳�� ��p��Z��/��D�{&}����H)'4��@�r���o-�=y��yW�d��/�Σ�%r�e��ЯzenZ��ɫh�ͺ��onA�L���Gh���~��'�eO��>���ۓ�]���$`�:�b�RK�ȹ�+���;��w}�06X.\p�2�`4vn�i1
:��_&�
���jN�\��1ʡ4�����o�r�k0F��G�O!"��uЮ�#\���8����ݩ���?�~��b��c#G~ei��Eʦ��� �$#�|2-��P��5�4���M��Bb{K 9��nW��|�[�$�hJd����d� k�������`����n�ve��C��i�,&����K�5΂�˲H#@?c[�4�G%Z��R=ZGI��ox�]󩈫������1hmXC���+��gY�j�%W�6�ǰz�C꛺Q�a�v��c��ǬJYhȗ>)�R�����V�*��xl���{���-��}{���=�`D�*��/��7�UF�kr��=�:��Wp��@�Cu��V��d0<1J�|F�u���6�\�.XT��а�N���?��1x;�W$�.dd�����aF��MjVn��u�L�8��ꗵ�V�D{�t�aݼ�ە���n��gv`����k/����xnV"�a�lÍx���y�&5������S�����r	����ѽ�l��z�
��J����.:�o*?­wbbu��&���e/�2c���{��.0�5_fy1\�3�2��ω����}����X��׊���΢���mw����Y�Cni��rwL�d�C(I^�PԷe�T!DQ�� n�ˢק�����ř�v�rٵ��x��=q�ڛx�j�n���)?���?@~�|����Ѵ�����g�͆�/���5�Zuw�Ϲ�0�!R�h���\#�l�.k�ɐ7��XCsʳr�K�-3+�;��Gⷌ��$bV�/��+���R��[>�1)uԬ�4b�2�7�Pq�?��ڦ�Q�C�[��g=Ҥ��2��;ĐD��D���9�K�>�`�[?�P � ᾘcH^宪�[H�<[2��Ct�B��p&�6Nt�t�
+�3z�X
�_�>d��r�g2sT��?��)�������bo(ȁW�1�M+s袆�3	���V�c��h5�qr	
5�V�u!����#Re>�<�O�.]��uc"Ů�x����L?bM�k�<��L�O����B�p�愀bw�u���,n	�{���D��^\\e������j�PI�F���e���:r_��9]"rq�A�>��v�ݽ,љG9� Nж�c��i<�m@�9Coꮷe���f �4�#C������#�����\������M�=�Dbo���1�+���� �Ӏ�޸Į�l
M��ި�ă�	�y�����Za��*�m��+����}.y��3�W�O��T��-�f�{`}YJ�:�k`z��&����	ԂM��	�ʸ�?_��#��|1W0�o!Ge�K�g�X�ETj��i�<��$j	\4��ס~�P�Tr<�<
�7}�w�jP=��à��^b��7���8Jpm�������}P��5���(��_D|�nQ�-�p�R�B+�J y9oc����E4��R�&(o���0K4���{<[�l5	��1��_�@��D��ā"h��2[lr(]���ɋ�J����<�����UK�T@I5ќ"�����!�	�p�\&8��AP
�^�Ӏ�d|�Z�1;ru�R�w�=�M�x�]�������/G��/8v�Y^ż���5I�o#��ńV�1�C��hW��I�a��������w����%����2.ۢa�+ 6��N4�s�M��_��M�f�8Bq���<��;D}���.o�i��"��<���������P�2�AnD{����ǣ;	��zb	��$Ai� �#�h�����x�H�_��p[��Q�=�m�/�UMCq���/��p��ٮ��T4��W��2y�bA�A.�{��S���u-��+yCk�Zq��Q�<�(�筞�%ha�Gv&�>j�g2yCG���և��k���kq$��X��;��������e@��O��ړ�~�&��1�qC�QT�5��H{R�:.�<A�.=��X�׭�jS��R�B!��7�2�0�	lB?�.׼�Qo�W��@o�Y'��/V�-I��:ȋ�Mћ�=d0Ⱥ�ە�*w^�.���<�}gY
3� ��O>�_�M+�~d�ì�(��r�0bo�#eL�� �G�C^VGr&}��k_�f4�,�A���D{�볊�7b$�'vǡ_Y��{9�ox�)���t�_}��OY�	kEG"}��)q�O�9Lq�_R�v�[��vd��j��Y�%�PbY���^N����ψ�_;wݸ�S���z2[(���%E�@W��	LE[c�c�|����|���Lʭmd0c���W���m$�sW�//C|�|�5��@+��yuQ���T}58����F�4k�7+t�aA�+�y��r�J��sX��>����Y�4���7t�ٶa.�'���Ք���֐��.��#�8����:��sa���hg\k]p�$�t�}�<�Y�N]�(
��G��4؆ݳ`s%UP�i��/6�q�*�E�MT.f]�Ӄ�u^�� �^�Ѩ�Y�\tTY^[@nKa�@�,Vϕڶ��J���ʲ��E��}R��t&���S �YSv�ĸ��f����A���wP<X��X��wY򌞕��8P�� DQ���k6��G�0��
�D����x���z��/�g�_�s��+��l×�
�C�R�cBsCI*��'?��t�U��w�ĉ(\������?����xr�$2f�@��c'-��"`XS�vP�uGy&S���;Sa��8O�Q�勰�q��5��;s�ް���	��0n���&��9���K��/�ټ��b�s�K�`�ç�����R2r�6�mf䒿�p�|���]�'p���J���%�B
�38k����U���}��-��h�Ez�|�J1@����s�f��} ��cۧ���o�)*8D�3�a���j���}���1|����P�
,H�%N�]���u�<�D����������t0Fȅ�P:�������/1�0֫O�0h#�#��Q�pĢ�Q��	y�I�8,��c�X:�3��שj]�nYa��-t��fHj�d^8 Q�D�����W��گ����`���VƠ�#`�.���l��x��bHW���P��8���9R����!�I���A:�v8�|�4r�9#$OEpnAk6 �?9��?�J�{�[6S���������j�$�ո�D;�D��K�/��v5���?1d5T��;M���v��AC����w��e3�$��O����J�)�h�U�K�b@��`^z�iwN9B�&	�x>K����2���k�D_�1�:4���М�#nX9,O9f������V��7%�K�CX�?�e���q�bV�L������,MH4�&0�s�x����`�"��F[\��i�9�9�vA�C���r+3t�q.j�(�.���G� 4��O�0��x˳vPd(���+2��������,�T�mv��(k��?Ȑ������}1�'����#��@�p,��@ly�k
d�ⓙ/[��:��3�������U'�\4jB��ѽh�߾4MF�~J(��=�@��U�}����z7j���_w�~�kU%k�KW�*/�.si(�p��D�����?<��qP�Zd����9��K�-��[A�6�С�JɆ�� ����&��B�q��UA����
5A���%\M+��^�$״����|(2��񠎏X&�-�_�5P�5vB�yڞ���D`�u1�����4��p/I�o�3�SxE��+��Ï���jL�����k3�bnrp&��q��SR���G����2@�K��]���{Rg�8����Fp��1�-�!�x�a��h��ln��i�tcjQ��"P.;ߋ�~@,��V���X���7ƿ�;Q�VY�����j��n"�g�>0L -c���Q�B���1�2;T }�����@����n>:a}U�F��a"��H���d�!�������"�6co邏���)��k ��y�2'�5�_������!�xhk}鲼UVr�b�e؋��7p���'���*���N��E� 'W����⏇R+Z����F}��tj_A�O��X	��D6���Y�G ij�^l��Tj�㭼cp�8���GM�I�I�~�%�q�ҮW�$�]<���]��� �U�C�~z��W���S�����H�r�צ��j���;���Ra�	�R	�v-\a�H
5���)'��,�F� �U�Hk�eC�4�@LUG�Ͽ���0wG�nŽi�Q��#��aߟԤ?M3c�=0A��]�V�,����s	�(�X����aq`��R<�C�Q�1#(���J�-��������^tM� g4��U�d�  _]�	@�^Ql~��
g]3��ѵ]b�����)4��21:�	���z�P>��6/F�P�Y��4v������J1�+YK��<�5�M,� ���@�E�C��㯘l�rG���C&5YI���:���rl`�+n��@�	�W�F��*���r��Z��˥u�
Z*��17u_Q����4���d��&H����zi��y�fQj�į�=-£'e��H�h ɹD(r�9�,S�]F��~ˣI@�Ӵ[���4��Da�~gU��4���2'�Ӯ�h�}/XJ∕��
�7��W3�G�(9إ�� 4.*C��������g�eLhQ���&���G��" ���G"u*�]����Z���P0\{��8�d޸��и���Q�v��J��a=�8��s��B��w�#�W��3J��E"�	9s;\�%7Gx��Tu�S�<�^J����§O�Um��؞���>W"�x8W��j~���Y��' p�j�!�	���]/`�ӡ=zr�	6�_TF3�觷��`DY�V4͝�`3�e������eH�f�$�Crl[�?J�����>�^�1�3�C��?���7���h:��*����E
O���U���{�4��=�5��~�N�x�����tʜm�1��J� d�n�p"�=I`�����������+�aY� ������ޱ�Q井��L�G�f<%-���q�M�:��Y.�d�ͦ&|����~K�ןh*�"�y��E.Y��Z��K�o%h��Ɍ��Ix��Ӭ�����R�n��b�Q�Ѻ(g�M�`W�+b����Ɍ�T�V���?��b�2)Ÿ'G^�o�ط{���;���Y�}���p��G�|$l�,�^�JK�X�k�Qk�ܫ�+I��K���P��1��&��n�\6EB�p�`���.k���y�	�>j5����n��+PC">�e�����9��Zg�~K���y�������{�,���iXtL��/�"�<����b�o�iG�#��}���._ˑ��SK8u�-6�k�]�;�e��n�?5�myw��!�g��a�ď�(~BE^ls�x��vݸ{!\�`� �x�$���M1
��tb��>���y���Jt���j��WFJb���DQ��鑨�\׶���S�M2hf�$n]�����Q��?u�Z���0�	��t����j$��J��⢖��6)c����X����#��'�72�3���Mހ)=��.��i��B�3�D�}�x8ċ��3Is�
��
Ğ���r��nQ��߹:�휠H���Ѣb�u�����G�1�S��h;�Ͽ�{�XE���%e �fD�lO��} ��HAF-��㱴f�� �.�\T� �5�`�L��`*�zM�b��n��n�X%,<j
,��*Dr��nC���ݸ�ZJ-��m#��VM!�h�p�@g#:B� �f����U��->�/y�b�?@u�$���GsH��L`Ɍ�����c�Rǖ�?���N�����;}�'��������U<UC��&��d~p���
�EAAѵ����_��Eq�˥�7������F��n�% �L��v��=��Tc��b��DM٧ã	o3Q�[�mo�>3�
�|�Gc�Yd/ƀ��RS9#9Ƒ?����y:�Y��SϾZ{:7���Vx#��d^�H]�T�n���ka�C8���6�r, �e���L�hx�M�g�Đ���� �u}��������D؎$�;�9�k�k@Rv����,N$��v������G�w�5�5>rjd����y���p6r$W�s!����x�Y��G���|
�U[ݓi��T4�w� ���S"��!�$�N_zY۠qq�4p��вǫV��PE�:���ނ�~����R�*��w�����r�~�ZO	$Q�~��'6~����y���GaRwwD ��Y�l���������޴�(�
/�z7�8��$`w�M`뗥'N�ӯ�Ho�O<iMQԬ��J}�U������D]�)�����MT/tɿ?��D��x����,,{����dЋr�Mĸ`�d����;�N^,=H��][�f5��x[�ރ8�(�#��>^�;�n'~�����3-�P����ͪcI���ќtˑ�{�Q��u8O��9��^��	�ٌq�tg�^_g���~��,j��Z�Kjk�ҥðW?�L���2�����~�=6,_���3�Nl[��� �a%/�h��M��Bj�-�Y\��VMI�>�Gb����Іm�BU8�ﾀ�S��r�xI�㲃 `N�\5��~�ߙ�v8�ٯ�.4Q�{�7=��?:i�N��{?r�\C�^-v���J</L'�L��}�������0���%	�R��S��nU�!�)}��M8Ք����KUv�.O��ߛm7��o�=��-�٢ղ;�L���2,��f�����TџLB�K��g�ٲ�u	��V�b�4 �ͧ��A8rX�9�@��i�J�s�]e�r���QBeeֈ���tt3M
ܩ/�PLm�f�w!b��Qd�fӦ{zz��q�̕㳠,�㨌�d!?3��8v.H[dŝ�`��4Ӿ���T5~�ɕm�ߔ+\rܢ����gy{^`�}_�B����.K�lz{���%���GsGa}!�֕��M�Q(Q���<���@����Yv�,�CCç��X�=��rc� �ɔ5%�~�5��k����u�t"���f��M��2��0����z��r��},P2S�Xlbv��n��:��H����)�8+�<C���@�����8,�ǁ--<�oW���>*�
%��� ��ǆ��[6���-��z��ɺk��)��1��3���)��R����[�S����Ş�f�m]�X�4U����9�Rf���d�"������RN�5�ϡ�ݷ��6�^"�V���:S��;�D�u5:��0���^�2��(wt{ý���L-�]�4�k��x'!ᵘ�U����W��o���^���~f��9���(�Zt�tz�.0d+8�.(�b���bʠ���!�0N�K!���v}�$o>^���ǳ������W����a߆��*�/���pܝ������M��ͫ�JR j�C� �̷ʓ>�j��\n�5ݛ��&��/�"��(�B�����^	���e�M|�`a!-[�W��-I�wD�������f�ը�BcO�<-x<[��(s8i
0&+���� "â>��>o.����\���q�I����J��;�C�/��S"yA��IcQa�����Z��S��N���=�u����j7]�������:�q+i���7�.�F���"ԇ�F<��>���xo�e�/?��\~j٨�`�%����g�{ͮ�L04�(�; ��������g)n'kC�ig}pY��t�l��%������p���k��1��x��ƟL�G���[(�:djk5�T�#���]����"��h�-�JK&~<[�m�I��&~A$]��[��`i=���.]\P����ۅ�%#8��'�iN����7�%�7����=���ΦvۂĞK[|/�u�(��}�&���zk'�s/���)��9��;v\��%kPկ	-<�hG�%J�c��YȀ}�x<�NA	��D�<�:��(�Ϋc�6�C�t��usz���8�:�peKO��e'�eJ�Y��)�m�٧P��th��4���sc��&���ˡl��`�<1���P�s�n��v/i1�بK�1���t��}���^�=a� ���C#6�v�>�O|0l��Ў�J��0������4���w�n��_ǡ2�y����ɤ�Do���� +Mi���VfH�0�����]`�T�:E�b9�t�0�P]��R1;��,�W�>�v֯�/�pwz��l?Z���\pD�*���(&p���L�;���4JU�Kц/�ݶ,����j��',��H�|ydhE�w�¸��Wl��
T�E�\���F�e��2�%X��4��3����l�>��� �f��E�^3�m)��\�S��f�=CDw��I�q�>/	Y�`Q��"��U��,��(QF���f�Y���G��Rl�}�����]G��ʤ��
"	[	.~�x>�!<�q�w��Ύc6�a ������d� ��p��1�e�!C T�W����A���ќq����w �;IU� c ��X֝�;[�%V%�V���_�o¦4�J����zSS~Gt�����+���D�;�+C�]\��]��k���U�Dl���/�h���G��p��e+�,�6�o���%]�|&�l�ؼ�	�)��X�
w��6�4Oq�<&t�Q����+-̰)�p���?�Y�L�3$���U!�IS�'�.�!�Bv|
0ze�
L/��K\kź���U4ˎ��X������T����*�4�Zt֥%�R���U��r�`�e��۽_j�"W�2���Ǆ�\ߝ>�:���E"����]DL�PWH�?�f'�A�r�+�,E#x�E��ہQ�����6�;o�emE�q�7���@�14&O %Lw��M�OO�g"��Y@k��҅���m]ȸh�W�'�1
fR	_k�Y
�Iǔ/��n��>ĭ$!d(��l�6~7y��rl����ӌY.���O��>i"��zU���>�۵��ǯB��U)aF3+Ƶ�s�P���R���7 f��N��g�óE�f��]܏�PHd��8�m�.u��ݚ�,}�s�MÈ��^4R0R�G�����TF�`�O{�'聝`�0�=��xE��;�7�f��q��+,*7T�D�j����F+�l�U�1Z�H;Z�(�૽�b�Ԫ���Sp��!��F|(�*j>?M�O����	*l
.������x�����̾�Ӗ��E���zL=U ���7�Cu�hI��Ğ��1�	�M�#)99d�wjЙ�k��!D[Rw` �����ڣ�+DJ�~L��,/dB���#�)�}E�,S�Q_D��ӀO��,�녾�4�`��'�m���z��z+�pG���V퍦+%0��y$�Z�m񚴋�����̜x�]��M��<K��ǔ��{��L93��&T!HV�����A������Q�{��	)$��0�O9��6_�ZKO���sY�.L������v�+�"�8p9�a.�rF��=�l,آ�����ŷ�,��W���(=�4��ÒM'����EZ:��!�����6��R�U�s��h���H�ow��'���c�nP� �%PIT����b#�=�gl-��H�|9}+�3h�	�E���2|���P��#��P�$�݌���,UH����À�m�G�˺�[��D�E��OK ㈺`4MX��:ΖcW�2�1�S�>h3�D�v�c0�1@�`w$�Z|!�zYa��.��]��pw��_��Ӝ��D^��\�l�f�.��A��^4�w-o���#G4p��1�-k�%Z�7TOs��x �
_Kjd� ��z�H��љ� ���Ż:�J�a�~j�%��j�������ib�ҫ
߄P%t5ҫr� �?\�F�gv�X�����0y>IXc��k����U�����s��xp2Z|=�n��40�n��㘿�Yp�*��d�#�������	�
vq��%����$�;��]{�_s��S�hoa�B���}��/�uYU:m���e�̎�5�R�'Ý�y����\�䬹fe���������;jb1(	ɦ���s���旝�."Y ����R!��g499"8θ7/mccL�K�g�O���Y���Y� EW�op5�n����楤�z����(7�$M|6��^mx�\����^ �Ռ��LS#?Z��H��@aFp��؏�����g��u_X�Qp���t�,)u�eV<��UC�s�k/(MU]*Ǧ+q���8����1!h@�=��/�)���pڗ��]�j�6�\<���.��u��}è�S_nψ�+%6��6H[�W��*H���ЕWL��5���y�7�&/A���%$'pF�V�˜y��M;�I"��ay�`���O��}y��h�EՐ����1�'�Y�}Lnτ7'���\1�O]�-ec[�� cKL>�]���3]Z��gN2x��������tj��h}��Q��q�i��Oz�������MJ^�'�7��>>�(a��[�v�����m��H�{������_IDDZO�����`	p�Â(;���;P�:����{�??�W�]���P[���u���z��1��$$1KA?O'ƺ�P]��'��B��<�*�` ��,�|.!g�7���$T�WZXhȌ�>���6��_U�.`k�0g�6���e2t���v���#*Cc���c2��A�W���
�(z1�l2R�+٧�� ����R���Lm͙��iy�e�5�5�� P��M�k��Sc��P+�cTM_T��r�s����L@�/���J�/�j�,�0Em�b�8��7��z1��Z_QG���F���v,�a���7����f>�|�C�I��3f���>{{$��Z�?�ɻ^�\"p�=��|4�Nd�Wz1�1��������#�ΕS�;�/�b9��3��X{h�a�+Ѵ�����>!d,�� �4��u��4q�%��q�cpl��k��Eo�m����+���$��/υ���|:.�:��w�_J�7����[\0�q�<\�4+ڡ���on�}�\ �nX�@
�F��}�G�&�u�ɒ����6`E�Q����>r`����6����Z���楦��O����]x���&�@`��)?ĵ��W��x��-L���MJ)�<���^W8�c}M0�X2F%�gI�#�޸ve����fpF����D��e2S���<�nN�������\��.�T����{"��E� ���Y<�u��S+��<�[%����kV�G�{�mh6`����]���r��Y7�V�d��~��ְ��
:D��FCvZ�������)�� ���fV�X�Ҷ[��i�U	�8`\���Z�S��b�^�Z���C5�X������77�%��|�I��,� �����lJ��co�*���>,1����H�w���z~P�k&/>_�wL(���2}{���ZO�FwA�9U%���N��{ZF��+��+�=��]ՙѺHH�����X�|L��
�8 	��4Mo5�ʯ,_���<�;��r�Gq�J0':�p5e�S��T���C��%d�E6I�~��@=��L�F��[e�ܺ��aǵ\�K��K�ܝdT�(��s�B���)�I,��z�<��9V.$c�ܲC�c'�ԓ�װ;#��J�@0~z�O.�E6��BD��p������ы[ϛ�V�(��7;%�P�ذ6�8ⴌq�@���M����gI��������
zč����zͬ��C�'U3W��:����.Y�	ʬ֥�o�h9��+��Hh,߉r��Fv>Ӈ2�,o�#��h�|K��1�"m?���vF�|g1�w�2�d`���;A�*ٶ�
�_��X�	���#&�I���{8��:@���Cg<��}�Z�ҹڴ�\}�^Ss<��x�w�bOE�W�����։@��j�
<Z��Q���K�+^�t��$ͨA�:�3���8W !���U�љ�G�Qɗ\����"�*�h��m���@\��'�/6�Y�#-��k�u-ᛀ+��pǮ�o�Ho�b�[V  ���ڸ�lECnU���>�U\�}�ב]�Y8�`�O
7��?(9{ �i�{_�������:�1e$J�a��*��b�o̕!f���ί��B|���Y�f�}��8V�'5",�K��?x����J���	�%��'Dr �����]�S_]���=E�s��u/��m������ �UZ,������|�0�V�=�:�ٔ��0���L�y����n�LX��F�����Icj����?�6N};�����a����n�(e<�է.�c9pS�Uܰ�زǏ�՛%��ލ��a�����R7�R��ʫ+4����)�UŴ/kj׼�gO�����B��K��-�y�7t����
.J��-N"3��2=��~�T��iwmH/W�t�A�̬�r��ΛT��C��sM<�)K�h�FV35L�X�q�b� DF�m�PL%8W��@L%��<�����&"��	[���[��}f"#=���W�_�?߷�^��a��.�27Vw��<�9��1&_��� A}���V{�A��a0}5d�[A��&8�/J�2�o1�����ћvl�wë�4����#ezM�:G�2Ȗ�hѫ��mY)'�7"q�4����&3��q�|�E��9 7��,��'�v�BR��c�b�i-x_�!qlΣ��\:_��t�?� ��B����\�������Q�6L�dC_L��h �Lt�0?n�	5�v��
���q�Ϗ-��J���s"`q�im"�g�5S/>0^_�b牲zf�����2�Y*�>.pE ]9d�Z.ߍE{F�#��y�m���9(��Gh}��Li�
�Q"f�oi�&:�ْ�X�(�����lA��~
�e�P���~�׏+�N8#*��4}�7�}�b��ϛҩ����MK~�t��fƗ���;�Tz�B_'�Ԏ�6�K	��"�����G��P�FƙT0��Y������~��+���@F^��o��&*9xk$�k�bi��&�sɳФ���U�*� Ć�(4>��?c�7�2-xr��/�-�b�pu/�Fkzp�46�F����G�ʑ�m��R"�!`*��~��z�0��/y�_l�S�'��r������c3F�n�߽�݇x���f�l�V]R ���	5�eu&������a蛾:�בO�E�('7�g�DCU�����&�n�!�Ԅ:��flr'e���ݫ�'�9Xj�,�c�4s��}�o��Kx�_�-d+ٺ��zcY��!_T�;����En�=���)���""��0�Y�Ѥ��&j !���+O���9:Jl�J� �f]J��s>���kl���­R������~F-;G�2�[ť㥫M�n"R'�j-y���4���;��`�K"Z%���P�PF!��>7��Z����L�����wAR�_\`2����2}f�4��+���E?"2Sj���Ob�'k��hU,��zL#�m��9�/��r��n��oʹ�b#��ʽ`҄�nKLhS��%&��(�5~����'W��!zg�E"ؒ����^�y	T�k<%Ñ�A���/S��{>Z�ͷ�Qs�fg�7��.�c�NBJp��J���~%z���=�VH��"��H�Д�t��`o���3`�գ�m>�P���dQ�3V\%g�61p�,���[䑵�r�ܔ�b$b���o[c�lsW�!zK�d�g�J{��DZ ���>GV�H�JJ,���wD���U��8��Z��"r��&����WO�x&=~��{�x���#8r�C�i�g´(�a��|����x*�%9"���G��i�yJq�`�j`аȨ�?]"�R�:�B�"���a�����'m�?W=��	ߏP�ܿ�W�k^�����Xp��O����l�D_:�F�^'�HB72f>��,�������[�y|�Q�O��ܒ��k:a�ew�sB���	�!8��8����$�a�B|y��H~�����0����Ou�q�������a�O��ɩ��ad����k?iѾ�p���Ŕ�r^-�á�� ���"���>F��qK�44�	\��R�2��iI�`>O1pM��Tos�o��s�yg됪�?�=�E���P��njvQT�2����w�SmAhd��\��:�,$�֦9^2/�A^�+��C�ү=���b����
�h:����6(w��Q��\(`�?�~�ʃ8�Ӽ�D\��!�
�{��^�>���#�qӝ�����ϳ��s�>�}Nԣ���%��֒���a	Uk�}=x)q�r
Y�쏩���X�ٝbd�n�g/>3'4����<V�W�6�k�(I����G����.Qi}D5e��gzU6����	��H5f_��B��T6.`n�d;���%�M �*�q�\|��(�9�l��wuܦ����9�/;���޷�x{��EX�K����?p�����Q-�R>X�jъѐ7�	��l���:M��d�(�}����s�*� NС�nsi��TG6��~PL*�̮ok�����[�
"��bQ����*��ΰ�}\�1��6t�{~�!���\�h'� �4[�M�4�l�3>W�D=�2���7	h[�˃����9�ZZ���m�A��O4gd�3���\����wH�_����(m�#O�J7�b���p����EÐw��Z�-�BH`a����_D<ջ���ڠ]y�1���&�O�iGD������z�[He"QAQb��1gh?��h`�b��[�N������L�/��A�c�N�
�#�� /ۈ.>��ȴ��*�{+o0+E`��&�����c����}qB̠�}������*����sn�����&�!���ѤҀ(�dp�:�u��dHi�SY*�O�^s%�y����]�:)9;Sw8U�d2�TC� ����$�.�-�6+Ӆ�I�	ئ���S�F6�N�6RW88B}Ņ��������8�.6�{%p�2&��Z�-A�G�S~b���A�4"�Ǫ�?Q��҈v-Wj����p��&����Tb�(���w�\=�M�j*�c�n�����`��p3����ߞ��&��F[f5!�i�DDezg���05�w6�,�����XO-�xp֪o��<�Y���#gE��)�*5���I^fuƓ炮¥�黿_S��&F>ȕG��4��Ȃ���)ɯ��+^*�:&P�%@���B�4��	������13����Rk��m�*���s֯2��\������O�:��y� �G�I�j��K~+¾�t/�p�?�:X�o��u�>���n�$P�uC�H�p��,a �ĥ/�[+I�����!��>c��ެz��|��������eQX
�A7l�J�@��	�^y�s�����){ii��pA�}XѪ3P���l[��ԬH��6�ڌ����t譇��Zi�M㺻$F1�F��U��)�dUw�?��c-%��m�(Y���c���G(�6�
�0q�@�f���]y;�.�u�f�z-@z}�++Ov/ĸ4�E�m	�8�QAx"�*��9d���d�d�Fiʾ�{5�ZiB>g��K�Q/U���Ǜ�<�Ǣ�y���09��&���˿]������(��� h��ap��;n�^�
ګ2:�����#,�<X^�����-��9k
 1;�;2��=ٗDc�i�wW�����KK��]e�с-j3������G���R7b���:���f�ҕ�D!=�OrJ�hȨ���	de��_����t����b��q���6���'�a�t�l-�6�;���ݍ���k3E䟀��סm�QP�Ӟ�TRWݾ&v-�"�.�T�E�ς<uNE-N\`���-!៺%���u�	��2��0Ɗ�noɫ"�Xv�`�����ՖL�����O^�_d�ʴ��޳��'������u��LwF������RL�V�S.��3Z��6dQrv�����}����$� d��6/�u��UC�.~����<\8�vʞ���t�����7����g)���ų��G�v��e��*]5^��ߢw�<V�
��&�w�H��U�!�n����=ʨ�b�}b�����X��oEL�=��=��k��e�Ta71�|g�H穡������v���d����_���AQ�Fq�"/=�e8Er��h����D̓��?D_��A_��`����!�5��`�Vc�xm:p ��Ъ~Q�R�ݠ��D�|�o~b�+X���RL�m����J,4�e�L$�J}�{�����Y+��m(Rr��j� �"�B3;����i���;i	���{`�7;:��N���W�#lV��`#Y�5x��`�M�~�\�9�7Ӈ 1 '�PF���1���^񅄷�:��!p�J҇���3��ì�J�	�C@�KM-�rx����3�:������:d�|5��o��=S�\�"�����K�T`�qV� 0a;|����S5�*Fal`ߙb���[�?��#���)���v�ُ�N����G�ch_Sy%��K�{�_��?�iܰK�O�H�f��n�U��oݝ莫��je�V3��qoN�x)k�S��xSه��(p�μ*~sՆ8',�*�����GѴh!jƐ�w�%�8β^� ��LP���5D�'G�Wjhc�����l�W��Ԍ�-���I��S���Un#(t��'͔���Q�F���u��5([ƀ�*�i��u����Q0ŝ#�GY�]>R��(HW0�p��d�Y��d��aڪ29΀c�k�n���:����d�P�,[�9= S*�^W���,'��7�z���⨗xd���E�㒑��)��J�
?Md�&����-wqRё=i�Z��媕����EfP�Qm �8��:^�),���X���yRq$V��]��������UT��&a<}�.$��hl�N�]AO`
m[&ы�Fչ�}/ڳ%�YJ�}p���6o&B���[_̕����|���Y٫�p���϶�I%w@^�f���𡂄��tz�Z~;*<筻�~�� �σ�Q����O�e
o��氦Ks	���Qj��j��h���Ȕ=E�b��S����d+��+�����b}��H7O�4����%9�q�?����!.���☓9V�Y*���]�����b��6a�T1�7�MM̅��2]��8&+u8 +rw��W��Tz;������훴&�H�9�����uz	�Lo�D�����'�֚O����6a=�ڸf�h�j�B�h���-z�:��_�?��Ha9$n�7�#�c(>2�W��AH9�|���f�9k�T�c��x�x#Ո��,r!�~�.�r��&�F7� �y��X����b����H���f{�g:���0B�$�O�qR�f
�b/����-�jh�akk��-���Z)�� �����䚏Ի�Z�E_�b�2k���&h�,2����l�R\�c�Qg��&/N�n�3q���T�Ũy�]�-6d�I�AF��� mT7�L����^�� �I֯|ك��J7���d`j����gV�g�%���cs]��B�
���r��J�i��:Ŷ�|���EO ��Xg�y�-���@)Q�O}��T(�{�(�{���E{@&V �H8
X��q�7�Y�����m����k1�tOY]��, ��JW�^4k��G��jk�OH&��I���Z�t��n��z��4!��-�����I�Y,n�Y���^�c�N�� Ģ+E�"=�!B�n�O����T�i<�
�(�X�|S�p{����%�a��z��/�3���S�y�I�$��J�ƺ�Ƌ(핷qcOWpo(���)WeB�!����@�`��,(�;� �(!��IW��Lqlm�dh?E^�����^_Ԟ��+�����w\�:�UĮ�+�A�f��{��\�H�����4:�b&Х��n�Q
�b=���R�k��a����{2! ]���]�?5�w�`��^$�����h4$�o��Kƣa��z ҹv��L������\q�|�Gn��*6���-y)�o�4���S2��H�F,��6ܒ�yL�<V[@�њrK
�g_.�G�F�e�?�,��0S������ܶ�2c�����g�}Al9M@��Pq����XS�x�e�����S��f4	5\f�����[9����#2}���\iw�A��ec{A:VD���.K���#'�2�N��*�������E�~B]�`�:Bl�*}_��=���������vv�͙6,��S����6h@+����w�qL�m-t����%����u1R4奨>��/T�4S��ʑ�U�h��9�#� ��7�xm�lc>����(�ǪmR.>���XL�^��[�J]2����xk��}(Ǟ�\;�}����Z-��{��<��}��� �R�l��u����9�e�.vB՚�T,9mh�h��h��2
���2����puh�,��Ujq�@9�����m{������8�n�{��6Q�W�$��;�Dr6-���җP'��C��Ʊ���ծQ-!� Pn���B�4׊��B�Eb�=����+�Z�B���\�~k��ĸH��D�>��J��nѻsG�T��6��W�O��8UP �����"�_"A2�n��װ�/^�:��%9`�s�W�-x��]\�9ǢP��*||/��6�9?%�Mv@K7ֱC��q.��O�y���2+�`�iGAh6{�\��)n��,������:\����Bf7�q���y?����3�����Y6�I�Kd�sft�y�����:;���FQ��<�8������/���<�*\�j���}�2倈u"�c���Nm�Noͷ �6J��n��b��O�~G�μÑ�~> �gJUw�$����	���o4��B�Xd[h���M̸�/"����~������^�
f�澶�v|�p
���U���*hŮ�B�\u+9��1U�TUi�bp��[���������X��[�v"-�idq�v�G���S/�*g)�I�[����Ƀ�:3�4�5i]��zܗ�u�xg��2~Z�9����z]/�Y.9|��&��)�A3�cV�(,cX ��L�w���s_9��&C�U�\� �y;u1
�sw�u�-(��]��b�d7�w�s�v��ǟ�'�ʛ�j�A��6N(W����$ ��xP�E^��Ѳ�n�	�pi����qR�+��`XXV��|a�[fC��x����"U�l�)V`�L�y�5k�B?M)���zT5���Үuu7/~�wP˨QR���h��ØG	c�*\�n`Ĳ"s%�\	��5kg0�Lh���&pQ��Ȝ�y�mkb��(��B=�*��+�P�j?e�
�̦�����##��GV���={*\�4��:5�M�jP�ېQI��C�s�B-D��e8Y>@��U�pī��<c~��z;�§����rS�d����n9\�kej0��,�1FDn��o	�����/�*�Q��mNoV
�ێ�d f�ޖ7�Ky�bO��'���($-��+6��YΥ�N�}��׭�7{h�ɹ�ǔ���<l䭢��Cx�Ǡ,��A�{P?2i�����f�S�X��J��>�fe�ta�o�.|6�L�~̃kl� F�bf+�TC%�����[w������I����U4J�s]Jd��'$���8�����s�C,�B�^����ӂ�ZBg��.+�=�+��E>�
T�u���m gG����t�0lV��]��Z�2��=A�6�Ev[8Z|<96ԣ�ּLq� �����X�F�t��͉��jz��F��Q��K�O�tj �e$�4�3����'�^qT�Mp��v�^��:w�'�CF޹�e���]f����uC�?@��q���#(�����F�1�k�yD��>HV'l�xi�%}���2b�H�|��-�t�sX�A��_�_c�Ý���C���;��|�'PE���^q��H!��e�`[#�q��I��,-V��� ���5|1\Ǫ�~�)���J2�X 'RdUJ1r�&|i� �uf4-�E�-��ŎPz-[�cH����/��4�.C05bF�������P3������BsP���$��o�W늟<I/b<!�,#���,�H��l��b���5�ä�+�U8�`u0�Y�p&�Ӭ�bwFᛘ�Cd����_��?G��r���q�GNVl����pxZgA�`ê�,��`������=O��;?�שR�R�%_z�3�yWDRj����+��C$>	<��J��39mE�	�MIt.�)��6�B�Z�*)��T��=j�#T�X�)j��}b�J�yCc�������O��!�9�M�S�Ҏ���J���s��#�,bt�+�R)�@�ҧ����^%/�����]�7��`��	���I/��"�%Y�"beûzlE'�?��}U&�	/����ę-` �bF�N�t0�nY,��ħ��\{��x88A�w��R��<��O{d��3�Q�����G`�bZ���)`��\��6��Úr*F�C���9�Z'_����u�jdeŐ�q�DC�~�� ���!�q�O]�H�V�E�n~��5X�N��AE]��뀥��x?�X0g)�}	�:{Z'�pӼ�B�/�d�gx�L��d�n[ـ�R��s���:cGo���Ԏ߫�umQh�f�tz����������'��^�Y$��zdr���wS�0�1�u�[2JA�t��*i�1����Kڟ���ߟ� n�֨�}�$~ep��6��Qj��V�����/�l]���k�h�l$KL"%�[߈m��������Z���������$��9��׿�?��˷y�π�B���W+���dQx!�"�w���8TW /�B���8͍��x�[����7��N��f#q�NCZjM꼢����Z�
9KR�^>N�?y\y�,��/��H����S����.��5�E[T!I�ꯘ+��։E*3FM�M�(])��D�i;��]5G���5��Rd���CO1YT�m� T�p2}��hQ{-!���Y{^1�a"�����s�a���,�g����3x�4���g����}�]�l�m������#�Ex2o9uv��tيyh
n�&w�Ὂa���}<ȴ⊼n��)�~���e��<>�O�ց&J��Y�G���F4Z�����s�Z�/�T��9���M|����p���L�9��P�T7�s� ��9���;Qe5�r8���|��K���0�2ㄧ3�֎�%6b��o⺡���U�X�>s����g@t�S�Sս���Qlu�G5�ͱG��P>�;����*up"M\�����*��C�v��x�қ�)�,q��i�B	�ؐ���<\cN��yH�UR�
V�b�ۡ]�mǌ�aI݁�7!�����c"[��7y����p����^|�`�n	z�V �	p=T�M!�z��5Yn�(~� �w�g;��^����������:�� �.���G����з#ح��ƺ�\���Q�EC�)3��>wp����.��v���F;���O'X)�����A���L�E�C�E�����E=%VY�il�J@\�Z6�f��F�Ѣ�;��� ������|[���#]��k�^�9�M�ͺ��Z�7�x����z>x�\��3(H��;^������s1O�%���t�@�{�cH�N�� ٱ�[� rMJbG�F�$ˬ�lY&q���c��;-XG�C)�ÆG��a<��2�9�A�p��5B.��������g����Q��-��zax�����H���:��عjj2H
?۱�	�컡�vMJ��K׭Pi�\�̧K�l���R�N�h��2.1b ��:)��K� �v�D��`7�AyA�Jt�Yj���W�EPo��l�s6�2���Lqj7�"BH�k��Nl��U���v�E)�Kա���(g)�}͇�ѥ
N����~C*��F��A'�~=��=�RB `��u�YcE3��݋��� �A������:�YZ׸U�ݠ=c3�����J�pS�������g�k�}?���:�q&k|�����)"��~[���	�O�*�`3�rߛ�	[u��<k6Y�8�3	&s��=��Q7��h��J���0T�<K��pN���uu�'�m;0,x��.>䥫�3�	�j��H�l$g�����%s�ޡ'�-�Қ��(������򲳸���Y��2]�n�i ���dF�R���:*�6<�F�y��;!Gȿt
STC���G�kf�zЫ�w�K�atw�	b����0�.(�UD\Mg*UuIҡPDYV[7iǝ��V�k/D��j���N�[����Q���C�H3y��dkl��4`��gA��PW��<�q�	+�i?����^ǟ��y��b��F@�b�tn(vα���6Z��y	�"�gz�H�ڄ-����ӘE�I.:���u��p�aS|@� _gVZJH�\ᷴ9�����b6n�I�/Ƒ=�$�����1��6��1�w���#�BG��&F�BkCԖ�5wfD�i�\��c����>j|u�j����(YG?�ۿ�[¬~�WP`�V.����E��igM @�Y��%�u�zyO�6��%ᒨ�:w��z�z�9����8-�=��
���9��P4c��̍~��$����C�r��Mї2�p-f �ً1�$lCm�d���8��]qq$�7yX�vۋY���~�����b2�1��p�V{��i�L�j˪��k|�4��Ю#���l��P��[�N� ;R�ND3��6�lS��݉ݹ�Ɓ@T�z����8@���l�zZ�B~�#Fs��1Ƶ4����)Q%��`�@��FE�Ux\��4k$���c6l5>(xi@5�8�]�~v����J{�Of���hI��ɺM�Ńo^g�Y��S���"��jf^�o�w�������J��٦�"%����p?U$�[@�Ҿ+�����(�K�Ǯ=ֽ� �8){�a��F F����>��E5�S�4������R+���s�`^�w�\�-���	Fm�5bx��[X��:�af�ny�^ߐ���BR���t��Y!M�����מ$A��K' ���	!�ӽJB4���74�e,'���q�|׉��r��+����ǆ�'-f�e�7Z��'�qB}G�ֶ9�K�P�c�.�ߌ��Ak��txX�,�PGh�9��ؒ���VC�q�*Ҫty�]�ߢ�� �nĶ(i�y�ܣ-ȫ�ao�r��S�&���s������F�Η�ca� �z�����{v�rk�I� [�����ʒH��Ӏހ���J�v��A�/�ܿ(w�ak�8��+S۴̖��-x��$��25�7�.�*�\v4C��/�g�Y�x�!�4���z��*�b*��cN蝖�ag.V�Tb0�(vR�ggu|���Ĥ��uoXׯP�:S�I�.�As�H�_��B3PJ���@� n�ficB�iP�mS��֫������O���k}.�z���<��/ ?�����]�����\S��;-��'"$�g��J�7=��Ҷ����=Xh��S?H���4���3U)�ղ�4���B�2�3��'�|8�<`��'S���4�/^��s�4Z_���K"xWV���6_�ah�Of�1�D�$v���E��9�w:�t�)�w!s�N�Ka=�h�1�%���h� ?�7�%�}-�nf��H�Q��Ź� =xh��F���q7�Tʧc��5�y�-�����κ
 ʈ�����)H��5��׀��S�E2�32w�&V���T��8�E�~�K������9��Uf�5y w�4�XI�/'Tb�6�mh�OA%H"e��V"��"��U�/>rH�޼]�cݗ'i«�M���=*�>�¼+�g� 5/��J�N"<��%���}$��&x�O7$T��[�]����R{dݦ\�}"��W:����!��/R�Y��%��KB���M���^��#��
1L�m
.�)Zz�WvR�%��]�1 �3i_#���J>�|R*{�N���F��1?�gi=L��=�6�[(Z1]75F���L���Y���㊩bQ����Ui 
���	�p���{B�������-�t@��|w�.�05r5B.��ɐ�����ƾ���PN5�:A��H*4��`W�`6�GT�m�m4��,���y)�H4�T\�$`���M4����ؠ�f[}�L8G%�3�a�k%�:i���J�B��G��i�P���D�sB�5gK5Q��w���p�k۱yxR�5���B�	�t�9���p�0��M�0"���`t�)1�'{~��y���q�b�i�8/nf൭��Մ�����mej[���!t)��'$�;3� �����ڒp�Ň��o��r-�Tk���F���vS�ܝA6t�$W_�Z����w����k�����It$}�_+6j"�V�\IӲ���P�Ҵ���qd-��q
�khŨeWC��S���C�t��|���$3P��H�R��g	���a�N݇�=U�g6d�/O���Oۆ,^��0���|�Ѫ�>�pW2�vJ�5�u�td���ض��|#aė:�p�L�x/e�	6�t���}n�D�����.��^{�ʶ�YdA=�o���/د#/dq�.6�G#��{E�\��e&�7NE����>�T,z�2�5�$[[#E�&���o0�'��dՎ�*�O^uq}�	a�k�d6���M�q���#��41�b���t�se^}6�&��o
J�¸�ĂV����1�1�LInH	)ײ�k��6�8���R�\��$dN�f %c.P�΋vAn���
��n�;�pm�_@D���~Юcj�٘�O����~a�E<Gڜ�o��!Gv>� \�W�w�I�}�+k��n+Ⱥ�b��4Dmq�(,�����,v����?��͙��?kz���r3+V3JF`L*�Wf�¼�P�-�U���QĂ�_�FQtZe�x�q����>��T�(��ȣ5��tr@�L]o[ΤA��DE��ɣ�-�������'��]�@�D�ˉku^�'�rג�cK}�����N7��vB����o�[ӵ��^]�'*�.%Q_3�� Ї��uE���WH� J�O8�ۜ(^s(z��6Mլ���S@*�l_��]�m#˹��	}�$�����kL�U�h��q�˔�tt>���Ӛԇ��2����jw��n�v�{	��x�0�Q^��SO�ܔ�|Z�lμ"�R֒�N���;CڂޓY
�I�I����'�Ծ���D�+�Q���;�tk��u�M�<�v9½4$�U�r�b�%x�)V���b���ڍF�&��"@��v�A�K�(=���t �&�篪���*���h]3W��H�q�¥� vG�Kȃ7%A�@_΂іv��+*p��)�ȑ��*�,eͰq�z_Q��y��o@��<�L1Z��V>R��7��(�k{e��wreR_����ڑ�=��]! �]!� Z�z3R�l�}�d��OS$��7[]��b��oԅc�2/ �/���O�/L���X����8�<��P�;������a�a��,��!�۩wPi ��V0ԉb� ��7V?|�@���/�<j��:�HyxC*�04r�Q�6 ���=�X�X$N,Gh�!ʱ�x��$���X����	qq e,�,k��/��@k�%�F��Y��07(z���]��lO�a��2�GNP�עZ`�t�:g:&�1��a�����i��e22������,����!�����?�<p{p6�1�	QEU��I�!�ҡ����qf�rq���(/=L�u6����,��m+�K�R�����+򸛢���赋�Oe�t���T���tXG$�9�ރ"Mu�̻����èz��Ӽ�K�q� ��1q*�O2m'L8������G�棹�~�Y�6?oM�c!B�HR��GC�0����w�8�M;A��\3;��C��1X�6��y�2&��`�Z�K��!�"п���]�7�u�$Ж�vIz�S<^�_(Q�>3n��f��4��Y;�b²�oT��-Mk�TDԾ�L
P��ze\+"(��e��w��ߗ������0G �b��c`�Ua(Z�[������I��e������#磃Ig�;AhIo����Nc�	W?Dg,Z&���#��s���a��^�Ѡ�(3���/�nU�^d�𹠵8m=W���E�qN�ݲ���h�����s�rBYw28}۵�p_�GVq�ڰ�GS�W[ 
�i+0i{Y�� �U�qX(ϔ���:�g�
�א�+��5U������;��>����|�'Jd-Pop���a�us���Z�u��n;K6�o��<�eB ��`d���܅��A�=[!Z� �!��k ����-�QO�!����q��P�'��dP��QQU��ש^��P1�@���*�*����
�>���˱�g�^gХ 3*��L�e����L�[�SgD��~�^���y?<�Atz3�G�m.�f�Ցe>�v�c���1$���vm���z��fӻ5*DH�U��U�֋U�-Ybep����qI�Ve�V��w����ca��4�}!�k��1K�(���:������L��B��-N��(C��-��,],He�s��0�����ԇ��k���(~J���z�����#�I�lw�M!�]m��s�!Yz@ͪ�r�N.,拲D1�Z\�~�����cB�F���}Ό�ٟ��5M"��^䅍���$�6�Y�#U�s:)rnYƸ��yvK�AG��p��an�K��]�O��{)ŀ-_���c�7U*׆�rn�
3����6�%y��6��G���A@��(��$&�R� g�T��5�>Q�` *��9�y5��޸ؗ��D}Ѱ�$��?<�LWq)��k �D�s�-�����MJ!�Nz�"�C���^5�X4��dp9CuiT��ʫ]��V%���%�|8�}7L�ӣ϶P�oD�T�S^`�@
9I?}φ��o��W�p��K'pz�Bf\Z��U=�X�@� ���c�F����R_Gr�l� �<��\���W�0�Q�~��I��(��W��)�0o~bLt�L�^3M6�� ��'v�_!|����^��R����3�*�.��Ш���K�d���+�YG[vX��������t�x�bs���=���:��$m5%_�yao���KF�ah�W�qiYq)D��	��4i�_����pE*�NB)4�������h��g �@���5�_s*���v����fֽM
�^���uY0ڦ^	����)�N/:Q���]I-[	�"?���{b����4�σg��x-0�I��e>�0x5�8�6Be��Hܷ�QY[���2S�(��H�r8yȼ��X{>(X���[��c��{���A��S�A�p�,�<��Ǜ6՚��\�pba���Č�D��D��I�!/�Z󟓆\X=��n�<\�Stt�K]!~j��L�K�����`5e0!*>����KÉ�AE�E�P�{�dDX0�!vخ�R�@@��=8�#T��?��<�j�}'�����Ar3�}'�k�ʖ7	 ��e��b쐭�rv��L�&_�m�mJa����֔o֙Z�DZ^�o%�� Vf	MO2�CR�sw�W����_����2n��:ݬDFqc>�$�$47��^��7%ˑse��TR��Too�%��������D�K�:0h�P��m���Qu!a��j��f�~�N榺za]�h�, �{�Ӄծ��rPX��gdҌb�Jǻb�5�x�Ioo΢
Yt�X����x�j����J�U+ɀ��-�rI����O4��z]�d�L,��i#+<ָ�E���/0�ҭ�g��A����T��������v����E�,|�Α(i�w������z%�9=���l�3"��/Mkh��o&E��I�)/��:�+�Q��e�D�0X�M��\�(C6���Z?��dq�vQ��z2�-�Hn1@���;'�=�MFf���-�䆅)�7�x��Qg�yf�E�4Ӱ�`�E��J��Y�gh% ��,g����P݇���7qz���g�Gc^ö�k�LG+� �L[ѫ���������e���զ�b�����g�����g��v�?Gʓf�s�P��]M[�].��[:."� H�E�'�(S'��'z.�L�<�̄h,��9E��B� 8��u4R���V��&�5^��k�Bz��šrȃ��m$"Ș������|��D�"m��e��8:���E�5���\��¤�&���b�q� Blג5�����_̠�Tģ�_���I�-?1L�7K=x���x�|�!�o��(��qw��Kh?M�_
SZ=�3�]��eTE&�Z��i3�v�$��=�`�*'R�����&�S2�^Kr �A�po���U��T,c�.��s�����
wX՘���\�b�$V���L�yR.}�=���,��Ppљ���9�e�%SC	���u��Ϯ��$r�e��H`a�ZF��ּ8�#X2�8��ɞ��E�U��Ƀ�TNSp�{�׌�π	sc��X �cPpT��T�@E���D�K!C�_>Fb�qQ�-#
j|1a��#k,3���	�p(�C���b�\c�~�����J��e�C�]Q�	d51P_���#F��W~�N��݆F�XJ��1]��/����5t��Q���2�5�.{�D�_i/�����	�u�T2�3�h^��f�pF�j����t�3!��A��� ���zQ���
*�%�׶��L��S[�x�y<��r�U�ƭ�s�a��ƶg�0̖T���#"�}�=Iz��6ɀ�;Y��(?�
�-��QBjaI�_�oO�m��1��4��� XcZ�C}�*�f��˽i|�%;�uHn	jO�׀�H@CK&\�_���N�R�y� b[1&i�w��c} R�_��d�D��߲���Zb��y:�ن��*��?uJ��2K�ל7��9�1vF߀0Q�z��� |H:'@�L6�/��S�@�����k����kBJ�c�}�u��2?w��VI0���gd����&�cT*YQ4�3	��U:'�|��[>����]]A��QQ����5���.mK͜��=W}���0�l��� q��BJg�}�ΐ�9BH`��z��Z�����RܐQ�B�k�J���	Ej�#��J)8��W�����M�~¿��o��^��`���M�y6p+�]z��w��{k�M��3�$b6����Gw]�� ��JIC�� S��S��Vc�"�C\�(u�.��å����(�,8�2}(s�l��Z2-�b��a��6���y��;D.SKǲÁ��[���-���B㾳L�0�-]�{�Q>�VCX�:TA���IE�C�P5��M��/eu�f�8������e,�n��p���[ᯥ�TO�X�$�������8 ��b��:�h���mʹɍD��� ����M&��<b<[ch�Vڪ6�$9^������+�M?�WE�ܪ��N� Z_���s��1'��N��N�/�c�.��N���?�) q�e�:�\�d�z�L���������x���Vc[o%�f1U}�Τ �}×޶:�Ri��pE�ʐǦQM�yV�i3�\�Xh� ���eK:�Ɖ,I�N�k`s_���=�J�L�}�������)���l�s�/H�J�]���lE�q�?��ܓ�~�|��"�F�����x�һ\VV+2�d�0���`���V\Wb5	9�}�c?�t\�d�J��G���ߏtu���r�+���-� l�i�;ݠ�s *�Y#�]�^?��t�ڪ߿�����]|����b�Ҽ��^l�E苃�`��I��9��왑��믂�e)\�C���.xg��M�^S�S��dK�7NVD4(�t��*��c^������Q�W���q�C2LjKwz��GI����HL������z�/��?4�=������#��TFϢ����^���]O^I�HMzX ��C�_!K� �k�/��(T�O���J���z� �����é�{1SvY�̟��(w��H���!�s��Ш�	�g�1�h��ۨ��.9;M=����T��kPt @�yUON������y⬘X�͑#��L�F��B��H���t��V�7"Cl�7i1�E��X����RQB�a�N�T=8��B�Q�tS�iw�s�v�S>(����������O�Hz��,,�~��bHF�9�X�>t�>�{�:ޤ��k7ρ�"X��(��f�+���9+9��W�\��?k�Z~x������>����U�[�݌l�QK�����C�����ah$�>��ݮ��0�C��1��]�V�Q�&�CMx�y
j^�������;g 7���^aǺާ2�6�{��|Ed�҄���/*���9���<E���e+��D���L�8�Z��B5Z�O���p_	��㙒�Ka�^q�bk�	8��-�Wa�8�=��D����_����z̬�Rd0q��W|������|�E���ZVv���I�$n,��Rz�������J�G��)Cٓ�0�A�T�|`��==�X�[ࡗĕu-�n�&Փ��������	3�
H!M����^5Ӛ���G�S��7j�Cr�^ؾ�؅T=nup�+s$؞ܪ��(�0�r���m��5iK�������ce�~u^�cDa��S�9�I&�,�6��{Rn��Q������ !'PEP��p��� _�����F4��~�&jXx���1�y[��fN��(�=$�UAJ�:G�p�af��,I��LxB ��_n�D�L�����d��l$ ���	;���ғ�<�rM),��ƪ�o�2з�6�,�Gj�����5�A4�m%��+��%��S�noҞ�5��w�u��+�O�����1U�ɻ^��QbN�{�!�1���(k��ool&׿���ȧ���cZ&����r�p&�#vͭ1LQ��P��L[����{
���g&齓�}6L�� �8� �*Y�8�{Joy0�ė4���z��/�����+�i[��.\2��J0�;&��v:@/��π�!��2�i�M�0�a�s�ƿ̨��>��	��sb{v�����ow��O���*)Y0?k_���N�jۦH������=�Ѻ���A:q4���;*U�]��	�0*E��φ����U��t�S�Y]��� �w�I>!��v#E�B{ճ�E�n�~ܖ���
��I���Ց��t&�]��s;MRՀ�,j_����U0��=Jp��4�5�2�|��-�?�B�?��L�@��E�Jj2��M5a\�Ԋ����B.����26�]nz��ވP�Q�쥁��H湒r!uc�>����א��tu}�j�^(��N C������}�!W���i���遻�����"�1D,g-�3���2r4W���i<@$+�a�b J�݉Q�����[E8�*�Q{�|}kWa.�p�[k_��U�q�2��k��f���e'K�D�2��9��[��G@����L��)/��t�lE>�?Z��{�e�b���(�Z�[�R6g�q�������3�+-j� &�z�a�h���h0R��~C\:�� v��� �@#V��C�7"%���N&��� �*U�G��(�����E�-��|a�ck�
���f�>K�5<���ri�7X�+/�֭�J�;ߧ�Q������M�où��qU���gH�=^Dh��K�8���'��S��ֵ�hl�kx4ӵ��hy4����&�n2�OОU6ڒ\~76�̅�y���<� �0�:lq��q�Ƭ��#��eG��� |�D��,�@���l����<.v=s]���w���FTکj�����C��w�E��3^B�����>b�kq�[�]!YZo�f&O�9�8t�pd��.g/��*d|B�E������F�I���Ve���Z��#hGoCw��e�%��oۍ MCL�3���l��Nt�^'R�{�v���nX@���U�m&���ߺ�oS�����m
�����Rt�7�͆q�my:u�1S�|��V�R��R���.8�9Iľ�J�	-#��n�]ؕW���dڹ�������Q4��^ Φ�K����x_޻��NZ{�`0�zTT�s�ψ��'k�E��'WȜ1+�7���%�s��!u���2s��D��.�� fD��S
mo�jNH�mNǫ	��Dϫ|�4z�p�t�@F_���]�,�n�u�><�ݞ�*a3�=-�J�E��̪2M
U�(�|�q�o,�0�I�����KX�MQ��a�ƿ� �:�N��z!�jF�Se�0\���_�;�}�a���fC�	��U���[p
�ܨz��;o8��	HϫnY-�#��F��s�ڰ�E��,��Q�?�V`�aR��~q�ظUV�X�4¸�%/�c�s󸕃Ƿ �%��H��-�KW���f�%�iݩ!�������@�,���&COC��<�C�n��sG��r9�<��#I��Y�.�am���c(�!K�

<��12�{ޭn
%��S1��p��]r ��"�;+m�R@z+گDf4*J�2�n�|��P3*){ۤ�E�c��6�L����,sb|Z�ɸ�k�n7K�+��e�<��+E��/�Hn*.1 ����Ods�a7�ߩ�*��h�,ݐ^����^�����>i�Tn�o�M)-�&I�S�{��l�
;��[H�yQc��7+��p"�.j��R�0p����)��?e�&���l�J�FB�	t�sVw-���c�w�E��P�~�ʕ�����RïƉ�p�r��5&o3�'��YX%v����=ydR:,�#UwjpT&��ǿ�(a��R���g2`�r(U�_�S�L�=�<)OJ!�i�L��SA-������P��,�69N"ͻ.A��iBzxց=��b`H�����{�KzZF���㞀ch���SP.��"���sv:l���}x"�y:������=m��fz�ɸ��'B��5���xp��Ho>�OwiJ�Z<
i�A{�$��!ߖ��*����H�a���5�H��v
~���8��y�|7>��2��V�<k褀r�9R��� ��[�'YE�N�I&D��5_�oY,ۛ�Q��nň�#{�����*jZ���i�E_��f0eS��$�m�n��7��%��^뽾�, �m�bv��d��Z�<������l���2����#��X��t��GF���!:�J��L"M���R/[�@r��f�����P����#���+�S�O����^�?�N+���R �1|�����|��i��a��!�cWk�	|���r��8~iF:+����ցL2����i�L�f[o������	�v�^�s�+g�ڎ�S�v0U�KKԓE��`5��g�͌*/q#ae�p�CA�^A]z[��P�� i*�\�%������jݎ*ͼ���}�u�آ�TW��1�3�G&9�7G6��
�L��N���9���~��!�CB���hW��P�c:̀�<KC��x��f�~�J/�.k1d�p���J��{���Q�;���b1]4�+�/^������j@�$�����B�����n���~1/ᯠ{����o+l>�Xa�(�K���m0ţ(���?:�FJeSt5�FT���䎗����?"F�Ȫup��f���=�����۾MϪN�y��[C<��V�i+4�y]uu��/۟(�������Ŗ�>��Qrfv}HF40H�َ݀�`��=j\M���˨P����V��壄�������<.�Fq5����^(F�����W��Qz�]�#[����ɻ>�)$Q���|q%+�
�H����A6��;v��P뇘��`�����<=%���`��4�"U�L		��j����bţ�z��,�lJH����'�n����(�lc��%5��+��y9y�2?OAѹ�����ye�b!5��ˬ��w�2�,�2AV�<��QR���U	l)���'��ũ�&�.�ڤ������m�A�����;���S�fb�������`t��;�W�����SׯP=&��MC2���{��y�]f�,��J�ƛl�FN���^���s��<Q�B�@�}J̉��|��Vj܋,�V0=����p��Z<�@]�jOjڒ�T3�%)W>l2)RQr'��B��#�ӟ�T���oa�rn�u���"�af]��ɗ���a�x"�������J�'#������&d����О�j_��kA�Б�D�s!�;iVd�{4�@o�4G��G��� 0j����?���ѽ���8��q�%|��Ɓr��f��#�820jok�����U�$�B��:�D��D;l��e���,4lgZʁ	�*I�]��`���0�k��Kft��dz�r�wA>T���]��24鯭=J�y3��NG�ov��_�舺ϱ��$���Xk)-��W�5�Ȼ�@��]}�f"�69����������q����KQ"�����%CK�����o�hK�>�.�{�4�U�&Ԡm�<6$�g٫-�O��`�J ?��22>x�+�#�Z̍�l�D,K-�Ԭ2kҭ���g�}���\vT��47<� y�j�~��K��dT&�Kw(=D>݀��\�� �e�G�D���?��	/^��7��GL;����@ψ!�U	��~�,�RS[q%�twٕ�M
���y�o��!�^�ck7.&��Dջ��f��&9�t�u��?���Fh��6���b�T����N��zeCGO<˂�
��Ᏹ�����-�i��~g���ɟ,�^*������N�"ڥY�nf��{tՇ�?�Wm�t�:K�L���WD0��R"�WF�+5���V o��ȱS�n%ݳd��f)Z~ʟ?4��\��Т�轷�����ϲ�!ԡ^��*GR9������=�N�h�6�Ky��I��u�X[t�0zvtZb8Z�#���zzaW��g�/k��6���Ou�.UX݀k�Ṡ#h6����} �Ŭ^���Wa`�]�0�n���fIP����i_��jۧ��=2Ո�HИZs��{$�Zĕ�!���T8<�_k%��<��=���Afg0^��b�pj�+aX���O_�QK��	I�1�*�h�>�r)����{�h�Bh.Ǌj��_�KB�*�&2���Bf3?�b8>:7��9D�u�/�|�����b���^-��\����6K�b�ݣ���@˲a�
K4�DI�.����ΞӍ��,���e{����KϩXjs����ΣD6��z�,���]U��YZ����@���Pn/{�e�0�V���-y��"�PSS�L�r�w�W9�5T<BŭU|�ւ��?/�����x�&*�3}�J�G� �O����t��`�a�|5-�i��J�O`]����6Ժm�M
��l`Rp�H�ӫ�]D�R�.��2�^ ���5k����[?.�9��$�)`�U��J8xG�P5��O[={Ͽ)8b�|� ���"����j��؍a�:�7��8%\�y3�+�S6��#�M���go1�T�-j�+������^�ǒ��DΞ�Y�Q�y���X���6;=��DW?|�J���H�s�Z�� $�o������q���~�� �"MRƫ�A.��W��&	���ٻqF�|e�� K���N�gj �ף��׺Z�fժ윶���W�VP�-ZH�*LK:p�����UEL��;#��ɬ���iS������}LЋJE�oVZ��Uuv�w���u�~���W@���f!AB.�D0�e)kY����r��LP@������ ��a���E���8+�ݮ�1ـ��}���9-
u�N�� B�j%���B�����`�Qek�s#W�q��g
q,]4�o�s{3�ä8#Bz�� �)p�MR��b۟Сa��TH��Qd9QV��g��MkL�p�J�� �s���jJ��S�FP>�1�"]��U����M t]L���<��g	d6��x�h>>��9'�J6���]�bjY�B��b�\ET���j�/�n�O�����	9"��XM̔k������:��&�fX��v�+k��k���.��X�q�
�t��c�+X|���K�)�L�ӵ��/���n�J�+n���}�^�j!�G"!�Ua�j����֜ҵY�o����,���z��B�dA��L�%��j�B�/|�%Ϝ�x�$�"+sls���s,��YqmI{S�l�'�ޞ�r������(�Bݷ��U��̭V\DB����y�T�����d���t����H�ql�LB�� �]L�N�hw%�xT$��g�u7�5|r��ZfJ�LT2�C�K�/��EcR��7��3���؇Lj�ʩ@by.6�lGC�O�of(�8]���Z�޹�R�v�j�o�$j�~h&R��gL���h�Yt���7��&I��p�� ������U��\=���L	�P�I��6A��`�����]�i�
ic/�0C6U�7��k�/��S�.\"���/؈�P�
 ���RH�ي(�^W��^�l^�@�N���vM,���}^KrV��COF�)�����H݋�Xx�掠��c�JE+>��zc|Ƭ�U�?��&�PX�l���-b���Q�Sͩ82Z>4�_���{��Ip��q�w���e��򉒲���[�[ƥ��}}A���ĳ{!���zxQs��P<;����8� ��d�2H��m����F~�V��Q���j�[�k�k��d���-Q�9#��j,-�cp��1X�H�M���!�"�W�L�g��`�]Z, ���`;eW]B��6eφ��6
���_�]����"��vN>|	��c������ɛ0݄�S�K� +L'����mh�~��2C(�Iy���0)����s�X���E�vK�I�����<��JMY�4���g����fU;�{S��HuƢ��sz�<J�޶i���ۇ�[IB���K��������B�h�����rG$K�~a�,Ȗ�^K9z}���b8K�� T0H8mip�!��2�� J�ꉥ4>�2`�1O���>���8���X7,�+�Vn��P����7��L+��`ۻE���z!g����kn��Iq�3�<����]eN�<X?=���yl�6�@5��p�0������90��o���2�{��;Y���{��R�Q��E����t	�N�X�DB��3F-�<3.��'?�S�dpɫ
iӾ�V�%Ly���������B͐bI������{���%��E-�ٶ�~�o�Z�#s&�><	߻ʎ��t��XjM��]��ᣭ%�
�K�Gh6�̒�������r4�U(���ij[�iې�е�X�=�bb�g�EK�2�"�2�
��O���������H���0�P龋�'^:���p�[��i�]�� M�����*� ��X橖a�,��� ت�/>�gp��P������K)��-�����bTH3a7�0�^T��iT&�_KH*Q_���xw�]�G�E���3s#�rR�|�)������\��[)&ݮJ;F��mX4�J²�ƾ=m�ʽ7Q7�3JmB�hNȵ_�×ˇ���Y�Z�*?,@�O�g6��Z��+��z���#M@h��_��2'�J���	����a5�����c[n!��tx��q.��N��6��)Ѻ����\��J!/��}�װ�A�dT���bl��]�׹���,��jV����OK:P�J���L����~���0�>�!tA��&�����%��cG�(h����ŦX���t��τ�����t���0���Z2Pu5O�-��<����m��Y�\㻡^�+m�M��u����������@j�,���k3(�!ۺ�4=������nN�N��]�yxw��]J
�0�$#Zln(D���]�n>�e��'� �x��3p�M�	h�s�`�*��Ī�7�m9fS���^�t@'�՟��eP��?�=�	�U`���kN�Y��Z���{���7����g��e,0���* ����s$�i|ȞK�r��1y`C:��C.�h��s���uq�a���  �\���p�cK��$̨o�]��C���B��n��b��&�(�	�Bu^Th�YAof���ב�I�x�A6��"�I�P��A�*B�/M�׸)���8h�[�jJ�ϧ2�	�F�[)e��G�p��{�=�e�h��1!2��8nn�|���-�#�T�)8������M�[e�����tߣ��\������[��yl�㲭���Z�m�Į����6ܠ���x�R������r3&�}.U�8�����W���c}��[DوY��č�.�����Y5�y��M^5io�.\A��Gs%�B��{����}s��Z�O�оA%�i��$�u��P/����w�/�z{�D,�L�K��s`�A��5�ˈ�<.�ɬ����<yX���;�b/��HD���,�Egơ�8QN�
��r	]�b�h�6d�)�B�����s J7=��gM#�>Ƴ�ݦ�@��V�S�[��_k=��}om�_���;n�X����YeU�Ǘl�z�28@<���4%mvM��&,�{�j��?;�����,��'� ��8�jS��x:���C�N����	J77,d.� #4�DPL��j�Y	W�~�cXm��ʮux2�+vk�����0f���˙��eh\q��������H��[(1�/����x�3�LYa�v��"F��X�&���[�W1o��=z@���*�����r1߻y(YW�X�=e��m��i9SL�x��=Şl2d������}�eo��){�x��=v�WE����^��߳��$�l��'iPO��@T��(���-+D�����wbd��"��X�XcZ��<��������*��}�n�=��5�3@������c\�}�W4%5�t��TPܝRS�Ba]���ʵ�g�0����@\��6&�>�����<χ���8�Z�i�~-����O龂!wt� ��o��p��k���ƅvf � ��X��:�<K�S�;��#�ce��eh{�y?o�����s����[�&2����rn+��[߲��V#���Pu�,��I�)�n ���yp,��
��.$!�w#,�Ⓡ�<���q%v����V\�T��i��3�d�̤[g��+��GU�Q�nÒ5���jN�^%�K:Y���^���i�J�bn��m�r(��|4U����V-�|71�	��r*q>�Y={�ܐ'���M>�r��ꦹX�����u�>ʿ�5j���	�YK�~�]hi1��aK�3?ԮT��jM��b%�R���:��o�$�
X�e�	���s�n!�\��5z�P~_�����4�����mE��þgd׺8�z��m؄�8�F굻,�I X �U;�!��]��>�+x�˫�RsD��^�N��db����ov>~3���S�ӎ�_�~��J�:��٥���/��C�k�-��c���N��#�B�1z���ѯz10�U�^<�o{b!��L����0�0�|��#�ۭk�!�c�t�C/�&~�@��8��&n���d�'�s�G�'��Auv '��t��\g9Zm-wd/�ؑ�ѱIă��\�g'���*T? #�Z�������zGu΀u�{�uoF](x�[�&�c�����D��N.�[�pQ���� ��fv���w3lnM>��\K���0�9��+gM<�%�D�ؿ֡Tl�&������"%Qu��DV�����..^J�Rګ�H!]P���rЧ-���W��,���5��N����e���D~����0���~��c���ō��E&/� ?�ҵ�Kd����6y]�~�bN�H|A\Y��^�ގs����yh/>��E%
�/�c�N�#��%}`;'��2��V�+�7-�Q/���ڱ?�ڿ�b�����<&���/$�س��K
(�r��mq�_��V��rT�K�Sr�
��i$�����i�
��0�I]��%C��O��ƫkJ���Ϊr>[KXH2�3�
fJ-��n��'��f8;�D?em#�l�棱\9� c[�:�x��*�nJ|�	jJ��Lr)�L#����!�th�sD*�u����L<(ox��A	n?FN��.���W��A�t8�iYxT��o}�.�
�	�L���[.g�fg��zq�3��Pջa��w�z#Oj\_���~=�t	*�o�M��D�)5w��Ň���gE"~��-t~�/������2���Y��4�X��
;xy1�z5Q,8.@�K�/��Z���Ac'�J��;ـ]����ph��'i�obp��ǆ!�&a�|C��6cH����Iĺ Q��!�O3���@>�A�f�2��b09�ȫ��Xs�4.�n���z�o�I�o�6������o׺�M
y��S�g%Pu��#�P%����͢L�jW>�zu]a������xS"�͝����-�?{O-"+�f�¡��aI��'�aY~��ˡY�'tԵ����
�]	��0=�%[��Z�����.pW�H��\�)��>��e�,D���W	P��%g���cc��@��2Z[Ɵv�}�bO��������+<��M+��`������uLg������60�p�x�R2����%�#�1����ɸ��lL�>	�tσ���v�^ك짼������@Hw��:4PB�`�@C�w0
��/�f[S_�����O�POr|+���ty��G9bm/l[J׻��[�᫯�;VD�J�-�B�7y���h n�k:Nq����8���Q�r���������9����0t��oG��u{��.vM�%�6�Kn�a����&�h�[��oՉ,=;
�&2����;2!/H�d���w�[pH������K�m�t�����B���$CE��+ݼO�NJj/���� !U)7�I�"֢�PH���ƨ($��>�?���Cx���ۢ�����Q�1Ma�w���lA�~W#�5��*1V2A��5���_n�`+�Yt�lhP�E�Zm"���:Zn-!>ՠ�B��d��B�BN:���ȭ#c���U$��ũ՜��Z��=&����R_�:�&�(�u�s��^�e�N3���:�>���WU�.rg׎��"U����������:�#D���U�� �,޼�|��4y��s��݈=	X��aT�#�W� Մ���n��*c,��2�'
t:��5�J�0IA�������ș�N�� (�O��uj�{�x���nJ,2��T���1�)ۚ�y�J��V�[�b N�e���j6���'��~�hy�:�k��n0be���D[��ա]zq�h׍^�yێB���Ճ�h�K��*����~#Z7Y�*�{݊�2�rTh��긛j��N]	q�ׅX�3��5=�r�[������l.����"�0]Cm2��d�|�9�.�b]A��z���x�w��2,��K���J����w`�8�)[3�xHF�"���AݒA�_N ��Kf^*�G<+����d��铞��XH��}�"�c"�u��X*�k^L]������_�5ȑ�	���B�F���ߚ"{û[�iA[(�OڹM*� ��p)�8��>Z��1E�q�;TV%�P�	ù	�֩]Fd������na�'d۾V�Ur/wo���b�i��>9�$d�>��^-I�ξaɊϊ��s`@�}.�U�:哐w�r�|��fG��f�2\]0o�$�*��Nc������D��.]eh���{K����]�\�tf=�Z�mmR��̨��1�6lV�uzMp ^�پ��<{IJ��Z�L � ,eJ<HF�
�q�E!��~7�S���[zs�PL�ZS�x�����ʕp�t��_�o�
ĢSg��M>)Jy��yOЃ��M�ef��œ�����>��o@%ΉC����@���4�~t��=�ݾ=����)+Nڠ�n�O�P�c���H_-_rA%�Qm���kc��U�FP����޳��)Y)� N���ޘ�\��)ώ�*���q7��N�0����4��*��hӯ��b{�<>�����b��-��Q�=p1�L�J/F5�#�v���Vv�1��J�g|̀��;� H�C��5=k�p6cj�w����~%��p��;6�PJz��o��K���[�S�5�z�#�̖��i!K��p�����[G�s�ܾ����13��/K��c�ܚc���(9ɿW����3��l[�z��(����ڱ�Au/�o���ͼ�����`�2�zW�4��Y���Y�غ�	 ��Q�2��tƶ�7����J�(
G��h�u��>Qȴ9)�_�<
��6R���.��%���،�W���p2���h�.�ǁ����?H��j�1�ΰ8`phl���z�ׄAj�>�@������C떺�O���=c���B��*@�F��#�/)���Äus9���@���c��2 l�Ao٪y��J�������1��9�����yέ���9�/��G���O/�HsK��X�2;7hr�_)�o&��q��~�SW��E��#�k�9!6�&�3�97��
��o��y��7G
`՗�4d8"һ��ڮo�j��B6=�^Z��{̧���B�+#�	�k1��6-�^H�6�ݲ�;��t �����H��퇂��?�O�х���\cf�Y"�r �^�X��|��<$92:�Ak�H+*[}3İ�����K����ޝ� wl��ղx/X# 8��[S<�I��A7�x�*,�l��2lL��=�.�7{4�.;*B��cׇ�ȷ��#<�:��t�`w�Ùf4�Sl���S�n��U�.�%M�Lt@o1�ψ*$�'���S8�����Ґ��`���'��S
1{\����)fW��Z��K�v��@0[ʦ+�|��>r��b��6AϜ�N�������'��Ȧӵ*�׎
K�+m:�#׷ŏ?�޽�/T�����IaN�y	��*x�@�	����Zk�mE��
�%�n
�q ͠~)}��N�[��X���v��u#."Ci�L��y�������]��u�k=�G�,��LpSn���"T���j��ђQ�����i����(�6:�%�����2����ĭ�º�g���w��	��ŉ(65+��{�(�ZN��{���(��B��&:�����Q�E��,�8���	��#M��ӯ�Z<����f(�bK^k��/�C߃?3[;��q	�V���%��Xh��^������/�&�e���R����\T\�B�����Mܝ2D�]��J�:�#ݔ¼V�NF�+�X���p|�X�
"�[����3*rj6�P��L
	��8��+��7�ё�#병�w�nR��4nw�X�oaJbT���� �ͧ%�@������bwC[��H�0���A;��J	hw�m1I1/��Оq�a�O!j�.��.^l�5U�"���&�ܵ�I]�^S'�n��h8'B�Xuz��~ZcKVմ J+ �<t���Etm�z�`���ҳ`�%�OU�4y�Sـss?�6Í[�*t�G\��-���U �B_���^!���+iGrx�R�5�fk���pd���tm�Y+X�=\�NFe/Fs�%e�+ʜ�s��Lc�p.��6V��u�d��(zS�k�ip��`������Lc��)�
)�R$�Crل7Z9��g]�ŏ�[/AV�����==Z�]c���$���[�M���R��݌.��W4Ի��5@�2�,�i�Rx��h�������x\aU�ތ�
�t���6���׋�$���?9fE�S8���cW�zw��~ڃ��ʡwp��2�{88[��GGP�_5��	��)���M&���Kl��� �u%�˒��,'��)g��6����t,��	���Y�?����m�����J��Є1y�A.5j���Sy黖�ރ l�i_�u���A~~��c�"��θJ	\�A|I'Na9��X6�sޡu�|¢�^b{q͎h�����}� �A��9L�Dn��H{�Et�؜�c�AuffK3膅Dad<8u15SV)?�b�ے�}���R�>��OiS�1��!p���oCm��KD�o���(?[�'������[>���zF��M>��;y�-��N�7�kI��>JN�k��J���FZ"y�����O ���!�#�n5j�*��ce7>0]��j��ϡ(��k��� ��s��g�v^L� ��@s�"Pw(@_�$�9D�3���+)鳋�N�R�L·��ZvKk�����/�@������)�a����"�q~l���[ؾNG��=:�N���Br�c�����F�����]�`��?�a�Z��H�h?p�-�P�F���9����'j��Kd"��]d��8Ld������9�R�hb>���w��6��~C�y�[o�,C�9_�,&�9)�'ԓa���R��R�ʟ[��e�m�\�EI*
g�'���1��%5�ꋑ�1�z�)#.?��)'{����j��(NC|P�^ ���fyJ�)�Q���
��el���0(+j����Ζ�*�AT�2RG�/���k!#��~�:p�{�˵f������S�pvq�!��(�Щ�Wő+�ۦ-�4{T�19�̊��Wu��#�d07D{*q�wл�d�ZW��/�q��K��y��̼��,���P?��ܻ�AA������T�N��3NꦵA@f�4��"$w���������mE(w��E�������إ�4 �TH�BP8�t��#��"�6 ���ұ�>q��8����~��;7@��Hb�� �g(r��Q9��pQ#��,��	�C��U�l
3?ՓB�<�^3o�v�ZgZ�� }�%�my��[���%0�Z	2�i��@��d�l(�0.�X7]��r�'ˠ؛s֠U�f���Pr�=4%�m������I/���7I��o�Ջ�%���=�Y��{�G�%QSN�P�+�y�R���"��[%$D]�n�������x{��r�89�O��a�~�R|NuI|��Z�YPN!5���fo�d�k�Lৣ=ô\tCo�9���2��(ѫʉ&FY���֐���Īi�D�פ㎕��x���zź��vx))�P��>UE!JI��� E�$��m�R@:�M$�1�`=����J���7�g�N�Ì(4R�M�����S�^s�z��b���n������B��f �e��_k@MA�4�hWO��:�F���(�,fTb�-SH:�cJHjS��x�&X`a����x�XzV9d������<^������B�<����<cH��OJ�e�4�U׭�ݸ�MiE���'�h�����:C� ��P��#�񑯡�@v��&%�re�SȐΠ/�_�S@
�&�<�h̓^����H��ͩ}��X�R;
ƌ������[�+�+�x��h�4��{	ɥ;�u�KNc��̕�<o����	�Ј�>��j�i}�;�y��г����\]_E�Q&G2U�=��bq,��Z�uR�q�`�c]��~�S�D��X�����!�\�X�xtS���\!a7�P�V���=���X��]�� :X��� ��&Wtpϭ.[��,֊|�,�����}L�o.�`��z��E���!_�oBx79��Ko��[�&t���խ���� 9t���)���@kƨ�*r���h|��d�7�Ul��`u:�Ęf�e��\B��Lm�_-t$�0}�xX�/x!��^�aBp�b�!b^^�}a6kD_hOD������ ���b/���z�3��u��Wf��C+��N ܥ�կw��ͯ�@/}���´�q��4���v�-���u�|GV�9�@{��)Dmj�S��彸�O9��T��
df�ϔ�D�/��8��)��κdk��'�IUi���B�xW���ev�ƭi,���Yzye���+JڊO���᧟�Q˹l���]}�C�(�)cw/�6n���#���MĈ f��qQ��@��������&}����웫��	DM���9�52�W�Q����屇J�u�qE��Rsg��kohF�0z��u���fY���<(�2��G�}^/�lG~{a����P�uη��:��2E����ڌQ���{�J] kÈ����t���X<8���G{��&؀�K��X�x��iAIp�(���Rk���1�A�*
J�3�>�a�S�nR�Z�;�{�U�K�B��-�W�ƽOc�/�ȽU*|�����̧��i�����5d�7���o���j	�������Eа���B�+�M�B($��Z&]��\�=��1��&��q3ܞ�^���ݵ7}�$Xs�L}��H�V��������jY����t���v0i�%)=LTɽ7��j�M�yK�>�:�%xB��q�$%�Y1�2!��+��<6����+�HָK�d%5q{T�	D"s2{z��4�usM�鱟Q�u3�{-Jn+��n�d�S���g%��[���'�N���D��]
60�_����F�["�d���l��{S��j�/����D��Mp��:0y�Ǟ�t��~W�Y�W�����GG������3N�E�����O\w�7��j�a�sn�BúL5�sy\�G�9NKwM�>l�l�kuH|s�����z,a1��#c�q{Ό��K�W�j>�u��)S���5iUj��uʣ�g]�f��V�Ԩ�x�����m��;┭r���fT÷���8��X��	�^Bm�ӧ��.��dA���L�A����Q��Ä�@��%/5h*wL���;P��%����FT�Ҋ��%	�{��삄$@���UB�ӭ:6zwK�|�z]�E����\:]j K���F� s�p�%�*G�U	�L��͕����_ϩ�֒�v�e��Z�[�t'��>���(��^G�暄-)���=���*VQ��ܸ�a��S9M(��#Ȼ 1����� $��;�J*|˺ /�Z8�2�[�]e7)I�'u5��-.h�ȼ�鄞$�LaS` bv�r+�N�&Şw�$Br3>�%�R�<ւɂs����Uc���.�̼���oض�d��9�&������H�=b��Z�:R.wh��m�[ߨ���k�1�=}��������#O�mN��� �e��L��m<U�qb�L��L����ͧ�.5���|p�x���4C�.㝁v�ۏo����J���կx%�0QJ��ȎR��UoBe�6����;�<Z<���6y���Щ�;��ks�pY��^������U��Z�d:��c��{�JƓ���=�q|�*
���6����c��#�QVE�n���X�����Ph�JH�����l�ۮ=��0=��"qN�{5<&�bxҫε���^���$�՝Xi���
��g=t������/�����d���1M"N��/��0�܅�c��'T;@���S���R�¸�LA,�х%�>(	_l����%x2��Z��ț�P� {#��#����܇�i��{��i�C�J��f�C�`(|g�޶;v��/�_�����A5�)9�v?{�回1�l˸��WU���(��%;s��Ȧ�c���Z$X�0o��-�Z����
"=�7�9T�H7�z!	��Ol0o�G��z^Dw��w�w�L�����6YZ}�nX��q��)(�+�&#9�]t�MY��!�K�l�P^:����a�ĻA�2[B��dI>溠��Y�I��B�&�t×��.Z*}���ƥ :h��3�^Oy�N���ѥ�����,=��y�Xj�:ʝ����!Қ$�������7u_&�f��沲���1k)��[�z�	 u�#��Njwi�b�<s ����-Ԫ_�R1��e�I���E]�/� ��1J�0h$���<)%��T@$H��_)�v[����F�h*��X�T����V��Ⓓz49yEsN�^nܦ%\�
����8���y�0$l���$�/�*p���ج��h����� �k��M'� �z��d���"����*
5��і��+]w\ñU1����Nꃙim�Fq��x+zZ�R�-��Q����=�.�0��Ge�4�|�5�('��ѵp��a=��V�S�bor?�nx�3����x�~�Т2��җGS�P�ǀ�!�75�\"��󭳈�4�%���8H��Y����OÐkU��ԊVұ��NEf'��[�֤��Ī��	k�C���j���e٩�sA�����0@87y�y�a��/��a�P�;2�ϚX����
o��5�Xy���ٹh��5���e�[����zml_��1х�޻��f/�~s>��b1*�l�v߫{��ג�QA@k����ay�}0���N`�2k�C]KK�Fk�$?w��N��/�W@yȜ��e��\����]�~�
m@��+��.3�c�< �!>�\�k3��`|^��`�' �� \���?o�f@�ǹt�g�)��8o�*��Qw�&��,BTQ�ߟ+��$�wwa�	z�$J)	WY˖2��s�blј�œ�O�U����C�t�`�s�F��5�ϩM��+52-{G� ���,V�}y�C|ù�չg`�i���S��?~�C��t�� �a��6�k܂|�s!BQs����3�H���x;̞-ʌ:Po3 HE<����x{%��(R8.�9����y���c^�w8U0:�ua�fRg��x��nQ=w�
&�4&��W��Ս��X>�c�m޻�1Ǣ�Anx�����A���1b����zU� �8&Mb��%�'���GD�B�2�u��~*�FfMk̇����(��I�������4v�#�b+v�s�	���=��r�C�7��D��t��X�"׶<%�b#�~L�di�����t����1]Y��z���
�ͽ��=@�d B��l�S�R��lOI'����N�Y�q�/�4����W�1����a3M�×�}݅=!+���E$a.�`RT�]��$[` }�In�����]��BlK=!�Y����h�
���7t����jZsR������?��?�Ҟ��S�Df�<�J�v�a��)m�Z���х�� ���Ծ[���/yi�Y��7p����o�)��̲39��rk�k��*U�X{Dco&���k�����8�K)��XO0���Sө���շG ��6=<_4�U���~��G���FT)��x��WpX�$���� H� �Q�~�{�����sZ�3"�$Yu"U]��:Ի�#enO�I��Y�:�hj?��%��`�����<`�d(s�\t5�'oEL����e!��1���6�`�;��g��4�^?��O���P�R=k1\$�8��͝�r\��y�2����):��e�\�N�ɐLqr�E95OL���n���U���&���~/�TH�����{}7�����+b@Æ^>-����Ծ `hA��g�~[M.�6�jZ�P��#�<���F�uμ�R�i�+��s�\3CD���Z�>-�-����Z��r�rB��+d'�N:(��G!�U�Z.�<S�e�&X�^���V�S\2yޒrc��B�}��-��I���Okj�{�9����ɺ�=���A��?ҳ�(�x�S�b/wq}$��+ގT���v���ɭ(��-�Pg.mL/������GH�؀a���חq,K����݌3��}�R1ScJ�c[PF�m��Ig�K�y��Xi9�u(�����rcդ�H�UA�C�U�vRR�d��{l�+	�k��
O�����k+�+\��0Ғ���Y��v1�1��-�I��^w�vȋ��Ϡ �5�\근k��q�d�/v7��m^�EB�C�ޔR�N��c��M)b߮�n+p��Ͽ+�>Ǚ]��֎�+���ѝ�=fIO�?p�t��@zX9�ȃ�X`��M���!G�����b�EY^��_���D��N�,�V Ƌ���]�蜵o����8
����R׺���[�5����eTEj���(��.2��ݪ�<�U͖p�lT{=��1�	(��Ou�|���:�>�cI���A�UZܱ�Ԝ�����)W	V�^P�}����.��>)�Up�����Z��ICt��w��e!S¯�^�@��obo:c���D(z����.�js�K*i(�C�t���/xi4m#4�[^����t��-�� �dj���R�=��1�n��ە+�+O�QZC���#7��( ߡ%j~*0��OZ(jpJm��演-�"}�"ϔ����l���QL�r�`�I�?�~�l��%�ر5c.\.�����lB�q�;���sZ�
�;@�'��b�F�](�k3û,pM����˄�s)_E���ˍ=���S�A��x�l+�/OL�\�E.�Д�'����~�����lN���>�?��!�qZ{�?�8�π�����[���2�\�W��6 {R�R�ҭ$�h��R����b�~;��l|51�NHF>�����5Mkll��n�d�k��4�;g<�T��t[E8-s�!L�$�* >xBV_,�1F��_TŞ_Ff�})�s4�N������}@��QN1���Ⱦ��4��� ���t���q�R��� G��7�cn�"�<W�@���ԣ�!a��K�:�I�<4@C=K����^{p%��᪨�ҚyeL?���+��m
2�N��u�>!t��}���:9�D�J-'+F�f*+����;t�Ra�&�]FD���<�J��+��f8��Č����;�-?d�O��G`���+��ѝ
Y��&}��	��c���oI�5�ࣔ�{^�q .WX�Ai�Ev\y̬�(=���(���[����|
Ym��~���_s9�F�5H/Xބ�w������J��ن��@(*ߵU���f�(�0��O� �i��x��W������u$"�ԱngF�s!�N2�,`�d0��p� �G���"zH'hwv����G��UTG�FwmzC�X!^=�Vy���G��q6����W<
j�����G�W�� S	�?�[i�g����� I=�»���]ƼK��>/�1���SyZ�����??̏������u bY.�Hhԣ#�}ĿLb���u����������O ~����E�N8���G0Mtl:� �,�	��k}P�̙͖y��'�����A������3.(m��쑚���h��ɔ��Vް��}��W�� 1�T�3-�Tʓv��ʂ���4!Cv�ິ��]�>��iG��.�J�9�/�>/`�JO%<q��({Z�GZo�i�3D���v3zY��:��/�T�^�y,v(!�r&^�i) j�E��I4�3�iK�E��0�:	= Q�b(���T"(�#�ܪ��PEGgL�(?��&�~-�#�֭����%��l*Ѓ�(�$<2<�%���<��zq
����VD'|��$��X�{�U9���/5&�+���$�y�'�i���nC$x ��SrbiY����d�Z��*/�+�4&t�b��)��l��K�G�@�/}k$��;�}>��+]�P=�<��Lx^,��lf����kY�	gU4ʵ���J3=���u�9����魸M���0��\��'�`�j������Q����|�N�� ��3�*�-J*#N�h[�_y�Õi&br�
��+ ��|���1�s���Ͽ
�{�r��3��^�y��a����"� ��N{8`[A!0zA�Ja�٧�_FoV��à��qf���(/f^w��C�e�m����ա��&t;�mOJ�-.�"n9W��M9���b�}.�+��� �x]+���39�+�[��boİI���l��W�B���`3�>��z�ZH{R48P��4�)�:�f��4D3ƨϹ'Q3u@��R��_�z�0��G�����c��`�Jf��g��.�"kK�&ӝ]�����tt����<
_�N��&( ��o�TC�0$�d1��NU]��*��)	|��nC�&1����1]��q������Ǿw�@��I�l�~��;�c�cZ�
=���ſ���-x�!��6D���̽KC�"�3TE���-��h8�����o�A��D:�M�t�2����7�b[�zE��n���4�a�o!�����N��9	=1U�H�������4�sM�s<d8�$��x���V2���=J��V�:������6ɷ��(�x9��PN3�:`��_������r���Mp����&�:;9[�ENm���𥤗���!�o�e@�_VR�F wf�����e��I��&{-^���)��ѥ�^䚽��󇋘�-i�ݧ{h�v���`q�|(_g�."Φ��n�M��{[[��|�:�t�B���nC��~BPѲL���}�*�R���D2����)J^��Z'�\�-~���zlB�{z�)���
�&؄��%�s������R�X��;a��uD�G��Sk*�ug	B	���Pǅ�:��nu����ĳ$K	�Yt��{4�\R��|���I�3�vfwun�hPx6�
M
�*LuRf����R8u/s#ӄz���̈́קQ �{v{Ay�;h<����Z��Q.\��Aʈ�|��,�F�;�;��g�����/�E�	��-�~=n�K:"O�B��~F"J�ky�]��bX
|b:04_�ɘ/�9�{�J�v?�ѣ�=��+� c��iZ\�4	���Nn/�������Rf������C�6[[+ȇ�kg�L쟕������+WD
����7����x�SԂ�!�&hɇ/� �cs/T{R#"7��yN/��)�ͮ�t(�tINd��a��Tp�a��ZJ��B3�Jǽ��N"�
T ˟?V?������&b�f���$�m9��ٿ?��bէ���#�������C�SH���g�6��#���k��=B�eo.��Ws#Ps��`���A�k��y�o���)��_C�����u�� hB�ǿ�S�-�'�F�Czl��fy�wx���ED��X����dO�큲�!���QmK2�٩�	�-��C>�#+�7��Gs�j��"s���-���'J��������ñ��nl1���di�?���0�������.��	0&P�6�mw ���k���M�Z��N^J�	����i�@�Z�����TX�8��+�Ջ�O��m�L����O�e*0��dWD�y3!���ˬ�&#�e�Dђ3� ����R�	�RI��JG���㬂'4�9��H��;t�4��-�\�*u�	�y���_��s�œA�y�^�8�`<U���>���
����nq��Ť뙦Ԗs8�`~O2���Z�*����߳Z)d9��dWM���(xU<�v�u="�)4����_|��gP9����p�*��-jW�銋9��� D��Q�C�k��N��gݘ���8j?���0�!!��@=��>!�h���Wu�K0���\��Ab\�ݽѴ��})�E:)�@��EϜL�r�P]t e?	2�8��ȏ��X<ܾ�}^�4����U"zT0*���|_�]n�����;0D�ρL�T���9���5���K��W��Ԁx@嚃��R����{O�{B�k�A���珟��I)�;�b��*�0m�m*bb��g����i�|�2s9r��#�u����k7>�~�/C����z����������\?�������x�M�s�� ���-|>,��#�Ҳ�;�b �Q�,'p �˼W
+ቡ��]~PHL�>�`�"�?��т�*-)�jF$�co���1\��Z�+>DBLw&�4���B-p.\�C'D4�V���;���+�@E"�?I���8��rDWn�-f�wʍ=��D{�׬:��<5$�q"��*�Qf�V�P�>ꛔcdH����#d�x����T%�8�J�B�8�jA��&Ŕ\�8�N�@��J��"gp=<]�x,�>�%�s�P�����7������Ӧ�VM���z&G#|dF��I:H�y��:��	��GhQ.�I|�W����F�P}/ǔ4����4<"�	����Xҍ�������x�r(���4�0�L��k����`O��F���9�.��S�ߔX����ƗY�US�O�G�����Wi�}����F*
4c�������]�ץH�f1H������Y�_d��� �K�⯹U��C���n�y�� ��g�H)e��[�v��OPS4.��H�d��u[�b��D�\�%ST��a*�)�T@bb�RZؔfZ��T�)�� ��{��~�T�[��n�j:�Zo���ǘ7)��{��HRj~	�< ���yޔ��{�ں]�=�N�!�6��g�����E.�6P$��>���0A�X��M.��?d��Ӈ���ZP���R�D̓H ��������h�?5�厰�pCj�Pд_�����J/q�dH���ܚ�����+�Ź�j#�[s@.0��[���>���	F�le�����ӝ���c�������T�Y!GԞ��WNԘ��p<�Gy�(�W�k�2n�(�C��/��kD��]�h�'�7��{���l!r�|GD�b�1���HhO:�9���Q��d�&�y\]ӻ��PZ�|�`��.&���r�}�<��ו�'a	s/���pMWp5����Ή�ۗ�_�E�ӡK�s0��p����&�w���]3z��'��ǿD7B�.H������%�,HoN��ФA�9�'�r�A�BN��a�{1g�!�n��ͺ�}��f`�׈�� �S5���G�ײ����bv�7��@���:�١�� �uwW�-5I*M-�r�R��T�������;d�JM�����;���9a����=�v����ngB�����=�e),/C���D?+��<���Rh[b�r8�`εAܲ����AFb��v�H#7�,S�9�:��/�si����g��zxD��K4��2TO��i[��a�;��i����{!T�1n�� ^�E�Ln�M��)�F��7Q�{�q&=��
>�ZՀ���;ޔCd�rQrLh����������g�{�U���pI1;2qn�b�lwa�����C�j��XN�Z��<n*��)��V���l�tg��0w9wT %L�j�z�l<&n@�d �ݟ,�-��@7�* �X�����ͦ�6Z�052,��`>��TvO�U80X8Y��\R���gsy:����˰C;�nR�-�Jp��5�SH�pב�<a,�	��v�D��<=�G=O_�Mn��%�B������|��g��K�40X�C,��V=� �,����<nB?a�O폎{7`��>�|!���4��3�}qW�E^��'�_Z�	_8��Q^���Ee�g�>�nETe�@a��؟��=�+V�ڟ��.���HG��7-�LHB����B䉁�<���[������o��.N�$'<RA��i7���B�T�y�����x*��gT����������}��)�KP�h�� b1;k�6��ǒ���\.
$#WC/�[��AN�~}��4���3.��n���a�A�ү��0q!��@3Q����-9s��z��������7�}���-�;�+O$M��E�_REB�SƩk����ǒ��{0\��H�}���wG�>��������F�n���ͻ��I�o�!���J�ʾEז���Lbf������c��4o��y�#��u������9�*�Oow9��wF����R[ʬ�g�a̆HD���0>J=.LQ �BjW+����c�HW�+�0���M�\}��郷CI�G¡�0(��刊�D��\���}�ҨgS[��/f%��l7�9�m�#/5���������.[����A<R��y*~zG9AE�I��$���z;��O�x�.���5{#�d��}E�.��]ܺ��9V�<'��8���l�k߽��UFγ�o�e�bgui���`�u㰸y�3�/��dݖ(QT�l5R�vO�h��N����Yw���o�bej�o6G�� 5��.������P��Jw�#YKHL4��|��F��c��	�ʹ���N]Q�ȋ`֟l)�G�O��6�=]
X���=iڝ��'{�j?]��@ԍ����j�$���h`����	H��io~�q��_}��D�Dׅ���v�O�K?�\��6'Y��" !xsS��b)N��p�-�#w#�.!�A�x˟Hr�>AIb����c���a* \0�Lǣ;L�����m��U����zU��kb${b���e�}��AF����d? FGͤ��Ϩ�Xc���p�"�|V��"xmCf�:_gH�5�f����2����J:�����4'QP_{[	�H�V+eoH��TffC�B�| ���T��=���(	�5����ԝ�<�Q&����hڌO'Ex�ё!���ؕ��!�v�ʺG�n�h\bE\_=�Ȥ�R�@��$!��4}��Y�c�{�<�3�0�=�u�T��5���8c�X�N<"N0��N�؄e����-�� �(+(��������"O3VƜ9s�!�g����؂����p;f�Vj�#}93��0�Ö�����w��_<�U�-�d�RfW7� ��hx$.�����ZZ�­ה!݉�{��柑�t��rt�����q�}v�PX��ߐ���&�l� O�y�������KL�.��0�i'���qX�$g�6G��g<P���H�/B�D �}lv��p��eJ�$	ܒ�	�a�zB�
�S3j9`���� )v�/��-�m�ɔʂe��]Y�_��!�*1���a?N�����<+!�%b)pհr�v�����tN��rWI�4Zx����Ȟ"���s��xˆ"����������'�ѝ_�(ګKmgܷ�'�Oh���8C����?�/؀j��P�V��
�?�]��"�>���4��B?��Z@7��M��}Øɗ^_���QQ�����)QYi�"�:P�0�tg7�3�Y^�pλ�:�"}8���y���\ӻ����6��ً2� י�n���-_$��%@X.roH�G�@�'��LDs��q	|[̠Tv��,��z�0@��T#?_I��u�GD�g�E�-�I�qF����� c��a4KWɒh1�� �hцʴ�ڛ�Y}'aᅣn���A�s���J�����q���'��a����y[8�M깸��I$���m��e%R*��d�в��[9\i��պr���@{��K<��}S�a�~>��feA��eⱘ�����Z���Z��e7�Qr��̠]���&������l?��a��	i�ih�M�[��!BB)a��"�X��HL/�F*Գ[OKYe�������;���� �'�?A�u�o����Fh�Q7�v��r�������9\C柈Z���0~
���$*6��6d��?�r��ǳ>�d�AA�)�=������"z�p���$��1=W�d%R+݀��2MVZ3�`����k �5��+%F������\u7����q+�0ΚO�Qu���⮞���#��ᨐ���r��c��=�K���R���ʉ�S�+8�,�2�wO1�問�(\����������vo�������M3���o�����K�;�aAh*�vQ FV�;1@���\�����&�
���� �S�m�&cUW5�Kh�2����"�t|�x�tW�v���.9���h	RAv:���
F��63c��by�m�(qϡU��/4N��I�1o�n�6s� s�LGj��� w� �JF��[���\�[�g��|������R<D���բ��1�Gê�f8=u�D�_1��U����jB�����*�
jٯ]��+d]&RnL���g�\�շ`��_�ϻ���txS�� �L�D�5�5ᤕU֙�}�y�Yf��9-�[��a
˄��.Y=���d�LVɴyYV�v���!ޮ�_AHD)W횎��˹���]���Mv�-m��>	�R�+v~��:���5q*_���,i,|��sx���ܷ���tq�v� J�Ľ�����'%�1C�*�M����Q5�`�FPt^RX�н纫��7�����S��_*'E�.����9���z?'�M~u�Η9Ĕ�/c;��W݌�;1� ߰-��L�X:��bcv~��>�ZkC�6k�ǃ"F��$t���/vih�D����[W���=K�'�?�*�̬,i�9t�w*-����cI��@T��Ɛ��5}�S������t�7̉,�!��0�;�g���"�^B�`�
֔aj��J���挏��L)I ��sU�n�d�~��f�rλ��r��C�6�Kie��s>�z�BF���F��F�4Ih�_�?C�x)J���Jݠ�ߴ�'�1�_���r ;hNR��z�H�q�O{��}N�*Q�_����!��	-Y��ˁ�g ^�!�xZ����{�� hT8���V�t!DN�f�����r��n���$Ó��0Ns0FWb�b�:4��%�	�Y�� �_��6㚓W�8 �cH�ת�����n�S��2�o=��X��C�ϱ�Ue�q~�n�y2���Pk�W�ݘq���+�L�i�T��h`�K7'�%Þ �a��|o���2m��O'�r�%����}M������vD�hR۶T�/*���!Q��Q���~ԹT�v�H)�җ7��<�a�W���M����q������7M��9}6�o�G
ED������OƷw+�zؑ\)����ATYҾ�E���4vM�L���q��x{���=JDj�����|�����Ҳ��8��� PlT���o_�t�,1��4��M�ʆn�����8\�Y��-/�jyg��qn���5t���
�O�TЏ<`sMY����6&�(b+:��P�F�y�8?��8<�[�L��Ϛ`����}~���W,s���?������ܟ.I��z;)Vw���-)�+?gC#����n,�G��x���*3�54JN������|(����&���]KK�-�pU�CBA�|?OrC��C9�H
�[H�A}R�
 ��ӐQ^<UU ��^��5�;��Y�^Y��JHo�� �i��v@�P4�����.�Y�"�O�yk�/��ވV�s�G��)k�eP�ƀ
�ê�{�D!��ؾj��7>�^ �8>\��t��������M,mkc1��h�ӊp�#�fm#=�����y�3"�B[�ck]W�T��$` 	蓕��ġ�O�i�N�LL�q���F�����3G~�|��k�_����<�۝���p(����`~��ߘ0�a��R�~�%�����s��MX���}�r��H:�����˴��#L �A��t T� ��<%}�s�,�߬�B\�?]�N��.݅%���{�`jM��/���8?����.����P�B�I�>�ޤ�5d�AC�F<���{y�զ���ƭ�6|�\9��M�l��)�&���R�⡑Q���wؽ��k�82\2f��m�<;STy%��E�s�XcBCG�FJ2�E˨���NeK�Z�|��[���L��g�w�$�m�8<戱R������R�z�]{�yC���7�X��i	5v�<=�#,�c�T2���#�H���X?S��_<���6���QDK��D�R��Ե�=:�u��F5���PB`8'̙'p�Xk#��\��2�M���T�_BN�rA)���� xl�����v��;��Z���s,��s���Gv��j&��Z�ۺ�RvS����f�wK�~|��&K�]Ⱦ���W����-����ad�AB��m�n<[��~��Ǔ"fjix� H�Bp_�I����K��>�?��D���-�t���K7 ����L�;^��<bn�`���s�����H07 ��b��%�tTd��s,�f�-F�?�Z�O�`\�̌0�w�G�����̕�n)�;���v�7n�53θ�����	[���'�����w��Յ��|�H���V�~.z��klgU���Z�Gݝ��<6��#P�6�a5�1-���%k܀R��ޙ���4��c���<���SW5��L8?��}e��n�]r��=�h1]=A�E�Xǯ�����ū�c��ɘk�|9�=o��tiQ�z-(���kK��Z�hr��n2��-y6��?����7����	'��v�+���⩎���r�q	�8?��ӏ|g�ҹ;����eR��hy�Z����F/sPm�ZZTd��f!�7OZ��@�Y��-���|B�L�e�I�,���2 ��z���(��^��l�6ƥG�y���� 6�:�<�΅#�/}�:C���v�Nk�7w������K�tw�+ѵ�N�5�귻o�ǭ��Z��s���U���V�z��ƨ0G���z3���վ7@@� �T/)��#3;�[VaL�s�!qz��5�5	c=��4�4�Xٞ�T�?4��T;�	I��QW��V��e�s�~�O��[��@�������&w\7�7}r�I&�g�$��_�:_�^�\J^�4���-}!Fd������w��l���y�%��'����u����=��Ԣ����I:M�5�� A��R]�R�Vw��h�9�p=6�d��n�\��T��M�^%	�$c���#�b�Da*&s��:89Zq��̇2T5`E,�s��� �ލ���jA���z?�O�W8%n��$���EPZ�m�t� #�-�;W����{p���0C�O��z���� -Ku8�@�%����w�xÜ�ü�����������8#:o�G��
��q���(Anr�_&V��u� Q�a����"T�Vi�|�k=8�w��,��<��h�Gz��I���j���@�e��蝰lM�QiI^�I;��#D����*Ņk�� )
<�9�	�Mⴴ��[���w{�א{��֐i�~m/b)Nȉ��P^�C�7�A04��?d�l�S��,E<�	��lb��S"���]5! RP��ұ��o/�Q�㖍���<V=1e���������I��5�Yy9Ho�Q��3������ZV��soqX��8�?f{WU���"C@�G�#l�/����dj n�A.j�?@�.l�~T����=Ǭ�F���b�N�(`"t�z��ͩ�H2{�S{!I�<�YI�o!"���@����Er@��T��(�t�Ns��	�fyρ.(���I��;�J�[�bt�>t}�4����	����4�X�pc:��ӸP0a����}gږ�✡Z=:���N`���J�����H�W�!k���i���=#�3�OʎY��k�D��p��q�s����\n���j�wT�
���RJ5`r�P��U���NP�`"�0���
��g�Dҗ���M������y4�y���
��6��4W�KYM���K��ŗg}��YW�L��7�G6ۓ,��2o�q���©>�F 4��df��N*a��?����0�Ӷ�&u�V����W�DI��s���,���l�@V�(��f2�_�ͮ4�g�<�-}����21��-Dk�rx����f��=�����,5�b��H��5�b�b��[�&�
D�B��؜�ES��hy
y�ҵ����v͋+'(����3�d��D��g��	O6c�ie��%���� �+k�����{n�	�*��	�S"ɺ�w�_Z�Ol��3/Z�d�"�+�]�:�V����2"sV+��&_0�k{������,�B�ul��4]�6|���-����7����Pb�:�O$��
dB�:���6��o X�T�S:�wS�J���iÉf�?y>�p"S.���6� Ix��v N���{�u$i)C7���:��Mi�Z3���';|C!7Y��A�O�-���5Tg����u��w��촦�`����5�i�<6<jZ��s�N��/Q�z�-�Ds���/j��&?��##;H#j`C ���R���l�d,MN-Xܖd�������w��a�y�?EL�b��L���~���_[�Mz'b��"7a�|��u�y��o��A��'���m�l�w��ݚYNqC�(,b�o�����녌U=�VFB{�6�A�zC���1A�S�������8rG��U&�$,�u�J���ԪW#H+�:�W��s��&!���p��!�T6L��I|��xe��N,7udb� dqO8�Dxڒ?\$ߡ�8i��(��+|����TW`�m�-+��*r��K��<�������W��>��Ѭ��$��9V��q_xq6�΍M����7����1�N����� �����F�Vw"��p�P7T�x�OÔ�C���E,�%��E�Sw�����㏃�'}Y+q=�ʛ��<�N�v�s�El"J9�j�Û�XH'1�H�C��D#��4�KH:��h���8�yʋF����ip�������!e�r�>J�TyU�\w�S��=�y�O	fV����,���s2�Ha�-F-V�5{]����oDq���a6I�{0ٕ>Yɤ���؊�/�lt��.�/Z*и~����n�6��
A�aJ�Kj'ir���3FU�ql���LT:{u�yVG�t�l���g�K���g���W�b��Br ��ǞʝŲ� ��"�ce�wC��½9"MDsc��愉��	/� �v����V�xkϘ���	)�-�;��������l�B�T���R������N%0Dm'�lvS	�jZl�@���$Zb1Ξ�uL�&�����A3y8S�c�|+	{�Ʀx����C-��U���hH�\�0n�WZ�(#�����cN����!����&��X��TIk�dy�P��	���8��0\���м�؅��t���E@�mpW>uy0�5����FBR�2?ES�6X��r��;��l��S���4�ښ��!���9�q0�Z���]{�3�˳Oo���-{<�.6_]�=X�wL�L �&��Y���*$����B;��䇋e�rCu��zHb�g��S��*�F�4/�1���d���!�ǃuC��
q.�_�r�>���>7Gd���FAW���_jW�����ɖ$1	 N�H�4�p"tTLGsҳ���f=�0��\�);L����ْ��gJ�"�]��7S�A"�%~�Z�7�2p�>�6+��m%0��n-�zjoL.)����i����/
�+\��+��ӞrI�
��F��T6�s����b�?y3���}#TR��eyZV@�LŰ�!y�J3�Q��\Y����D�da�ۓQ�L/
�������i�U��C��M�]��qt�� �{����E�%���TD�~��s�W�������l�L%�WT+B'�����5��+�i�l᾿�9���������ų�>�_S �/ğ�&D�1}捈q�_ޝS��.�?�~@keq1�=4�(���8�O��K	�a�qt���m*�ҕ�իf�@���^/G&T��b��ê��ț��C�-*L��<�r��Vj��q�D��w�i���U���t
�~n���������꾙+xQ�J�7X�`���:ĴQ ���G�1Ee/�E����q�'N����6<}sOM������@t��4=����^�+�]��/�9����Ub�էnJ	r�#�Q����yI�i�6��3�Zi�sY#f`��cMM[pg޹��@�M14�	��]��7���4gtdWR,|�qs0�@.���o:�Ha���6�KH���V;�pt�u��nJ�"x@:�-��n���Oe�ǭ�!�%���qm��*X�y�6��H;٥z8�K��&�[����d!ƣ�5�� ����lRZ"9����ظ���q3�0كd³{�A�"�BH��?�i�?2��g]n�/�k�x+̞�_�|��0����a��%��,�@��}1yN����\�5��~��0�o�#\ISB���P"u������,����K؁`t|�� �HM�J�|��ͯ=�7�ܞ �t �b���h��G�J^��������b����L�N٥��ְw ��9.���?^|W�x���'���� A�h�ym���q���:�n�g�p����������04XGW�7f�f�[�*q��xy�|զ�̜��$-=��FS�\���.�=���UY���+>�']ܑVG������
����oD��KɗT�`��D�S��u,��8���� �̈́gs���`I������w"�wz��uQ�)0�	pH�ߟ�m��蹻VW��p��F�^H��KU��K�[�0YUܐZۅ��9��J�#o����TEd�4,��&��{mD�EZo��k-�t�:3�(|�����������/w�*a�(:�;��-&{>�%��-O8r�����jv���Ɠ6�/T���Ϻ�����Ъ�"���=>*�e���atJ�֒Nw���C�"/m�Y�;�0tKLm�y��da"j���Ї�� :B6�l�l��0\&���<> �lR�L�rl�lZ/��1��&��O����^�N�|"�DǱ�l<;�ȓ��&�܈k"hu�� 8��u��N�j�mxʭC�{�Z������q��j~x7�z{D������@h��=!�e�*�d�ۢ��r�����}��T"�q�z�a�����MߍȈ�we����%,vA���^-��.}t��(!�g����S�f1����^��t�dJfO�W���J�BKb��u��O�k��n�л�"#�C��Ycκ��4ǔ*�ባ����W���A�I�"�7���FMf\6��=��	8�+I�2;���ȯn��R~�8��0�=Ove�=Y�D�e~��A��f)$\�icR����y����ܖ'i�<������/Ɖ�qR[�=^p���?L�*�LCQ7k���9���N�]U4s$(K�hb#�9t���efw3�l�%x���:��@�����UN	VAk�X��s\����4n=�k��'�ς�5�oq�*J��WS����l�l(
p\=��*�|��[�q,y�?Vc��ִ��>7����!m��$�Ѽ�c����R���_�=�?�
a4��͐P�*�kJ�AJ���te�Hء�Oq�Z}���`2�c��+�S��J�v��j��G��� ��i���F0 �f�m��ʈ����T�X�9��.����Ɋ-�d��W�iz��9%t�S�y��֔�#�T]� k��<��qV	L��wTS��g���j�������]w�K@��W�^'aEU�_sf^�MN2	?Gߍ�p~~��'Y���Ԡ����"\�諾���BS5��|}(1���*3�uiK�xU�3+�i;#����+�B���:�\F�כv�퐸<�|��"[�FJ�VIg-_Jsl7{�vK���[C �������>�u��I�j�n&
��/t3��9T�;hwk%�E�_��C8O��^���B�ۀ�ֆx�z�L�+��]䭝���;�܎�o��	��F�4^�>%�$�U/�
"Z��.�U'��]AR�u0������9���&�u_��a����u��Z[޿W�{֜��zl��Iv�����ʁ���H�����X9���s����?�� �1k�k.y:\�_!�'���W� �,�]}l<��l�|�LM��L�D��{� �gY���������,w�/
���u�͗u�����)�p�I	�� g+�T3q���0#v���������d�Ql,~*	�|k�c��q����G_x�`�j�?i �MV�-�¸��ϐ0c����s�w��d0�a�d֟���m��?0y�sVVc����.������In|H��y��j�=��>�;����풾�._4�:���VyQ%�S'o.3�ǘ��ݰޚ?��cA �Lސ���l���Q����1���<�o���)3��!Sl��Yx��
0Yb*�Lx/�tk/?1;�,���W�:FP�����U-���|�~x��U�P�T��	9I=�2�7�E�����l�C%0�y_D���a�S(1�+>F4V2�z�`��oK�u�P0�W�����/X4��-����1X��L-@O۠cw���gB旋J!�tP����^���'Z���E�hT$G�Gp���Ӂ1���ou�����ST'd��U�"_]|hj��3�	�æ暰������ߖ��r?��Ӛ.[2?vd����dC�ڕ
5K�s�dsE��w�3+���]C׳�ѡ�q�m~b+�B�?(��Q��B��3�������坁�cC��J'��}��G��c�$$�,4�Ћ�D�x#��8�����L ��A�i̤dT��' o�-8�]n�Qi�?Iz�v ��5�?o��QEh�Z- 
��]
�+��k0^��88w��LH�p:���~X'�mї�V
f[rD����b��5�X���x�����D���F�L��D��ӣ�7�F q�ZA�����5Zt{���{��)�ߙ��݋x7����=o9/�,zɱˁ��ЛB�S0M5;�2�6���i��f�~ȑ%��0�z��2�G[� c/��"��})? �ƽK�f7=V�e��^���iW��4E�[:�kn~\���0ׁa[�c%�-C�
:$Blh�����-6�hç.��p��g�����TDapH�u;=y�ktY������}�5i71d�D�ML����"��P�2���\�S��R���vyHh�9��42�0�����NH������g,s;ݪߕ�0q͵�~��k���h����0�4�)B����=��lӟ��(�Tf�&����m=mB���쵈=��n�Wt�H��1�T��a���Oo��DV��x$��Y�R�A}��iӨ����6r�!��:��ӛ��ЙRv148>�fj��RK��uԃ�P��a���F�'�1��BE����6(�u4I	۳2S�.�L��&V���gѻm�y�w��,��aF����u�ь�AE]��Z����ڮ:0�>�C�p�bF�`�HϮ��2�Vy�C���ێ&�Қ:���H�3,�u��U{�X�m�v <�rR{'qVU�����|DJn|�,}f o�dXKj�J�	Mem ��*0�ggP���v�d�e��~�6?z����h��#b�����~ck䰿�������
W��8_y��W�ŌV��b}����;����mg�A�S���҃/�����kܗ>V�Ҿv[E�/N�EY[���v2oS�Y3���B�uP���aX����G�W�๨|�"�d{̠G�Sԥ�Dn&�@P�'�P�k����RF�Aߊ�≲9C������q��௪}���*b]�8׀iUK˿��I�D)�Dǜ��获yS�X���2={)v҈K�u���D����D�y�-�B	�e��Qo'mx�L���i)1�����9��D��,����s�
UT��ӧ�?��,�j�q��{��	���|�~�QM�ޅ�&���%v�?�W�ic��PLUƉ���p��9V��<ث��]�*>}�w N4���	�1�G�ag�	\)�3 �.�g���2�$,.c�Vi����4S��q�ˮ{�58uph�jJW��c�~b��a��'S:��E0q�5ҩ����z��ޙT-rƿ
/�Z�R.�iwa�]!���1?_�4*ި).E/�M�Y�T��u�΂�xe����:��1l:�Ƥ��::�ڕ�O\��.8׎u��V5Ǻ�v$S��y�b�`�� Ok��?�;e�9{�\9D���Fl1�s*8�gp�n���yl
�'j�IML�᷸(��{v@MS)�SDf���܂��9��>'(��qpW�L8�v�ˈJ'2�X�v_X3#M��`����8�8k��T��#��<bB;�=���}���� �����g��Zm�yae3?�l�KrE-{-Zm���3E5�Y��k�0�a�L"������&x経�B�ћ�/�����@��\��\5s��2�&^!^���%��)��r�����d��J�S#H���.o,�$h���*g���hT*9uN=����̋'�Q�ј�Bm~#�O�;���jN�;K�)�p��ֲ��Z��_�����?$��j��:��]�&�`�TL�Fk��P_	a'�vT+%>���<Lk~�إ�%�
��l>�Pz5,ap^��K��!�F%��Z�W������I��d����l$�2;���̐��"�Z%&J�3o��!	���I�#�D�z� +kT���Q���ʻg��6�^%7��0�eJ���R��#t/��!{@)l�ڃ1tr;���O��G��Y+��Uw��Bg�ۓ�)z8��*�:5ӽ2����*�9mTC����".��NP��g��o#[5�<��/U�1��Վ�����o�o"���%�C���'� sS�>w^�f�ʩ}D�FQ��LSo�>�Zh������Q��ع��g�ꍋ9�������C7�K�b潔�s��ҧS
bv�;ex�� �$��h�ᄹ�k��֌�6����`��GM�����a��&\��ت��-�|�}��EqK����l)��TK�h	8�C��U��|pa�mw�>��+���_J?m����<��+Mᜳ�p,� �}��vs�rUi�/m�ss�����
�Y�A�D��#2"�A <岦VJ�Z��C�;�r��R����I����~�^��#��ڼ<����J��}hYׯx g� ^���P������/�϶�N���F���MZ����Vꚹ�a�S���1276�$�0o-vWRw)�����ƪL�1�h�z�����nIH�Ty.׭���q��8J�C	+�P����U�R����>�n<��\��n<I�o���h8.�s�D9���4W�t8�]�g&�c˫�B�T���?%Z{�9B�B�&/�@0����a��ێ�n��	�W��n"q{�d{=���x, �p�s,é�}4zz��M��G��\�-��80هh�,b.I&�KF΃xL���<�zcj4:�4j��n͚-<�?�`#��I7��5����5=�a[�5�E�	�D�u��r/�"����3�p���R-�h>��'�c��	.�
��ì�:�ƨ��  ��q��Ѕ_7�ZwZ��&����5��U6X�8`�u��M_���O
���[2��Fj���pZ醙�Q>a��?c\{�- ��9��ۢӲ�Th�'�C��7�\��/͖S���������+F-c�˩{��
��]����߯���Mff~�`���(Hk(i/iO�	�b)��g�X��T����>c0�?�X�5�lي',���}
��L��*c����;��mqҟ���,�rQ���	�<K8gg5ʁ��������D���e
z�)ZEj�b��c���!��o���{=��2�G�	C R�[��X�i�>(���|�[+���y��g%��Rv��u"�;o^�F������M�YxVA�՚���B��:����"�+l��{�x�P�yI���EKYo �Xļ��o��RF�0cy�hd�> ��7�L|��gV��Sr|$C�wX��so=��)ͺ�-&�?������Ł�x2]�J�	�`��.�$�����Xg��a�����l �Y� Z������J��_�R�3��@s<�dߎ��\�Q�F������w�?�M?���m:�|�N�1#��	Os�5�A�\'cQ������U���"��8��E�-hq�U��/um1�����Tg���_���&�cb���+~9̔��˸����K���b��lfD��Ӊ��قv<�,B&"��'5	���A�%�'U�,nZLϽ�G��4=b�-���!T(�cl�&��vQS:�O�g�P(����䘭�쳜Foڃ�3y��G8�f��V��5����VJ������L�-P��*��V��b���A����v�e��)���@5?��oy�=�mX���^���ԟ��OAj�	0}y�T�3C��������J��X���6����ڈu<���j��y����`J�o�6�F��e��M��%����.=�\5C�Ω��=�-�R6K�@� ��WoX����ɯ]�N�\�����C����J&��#k�R$������>F��?���{�U�c�V�>HN+�
�o�VH$�~�.����s>l�����o�.�bI��7��v1M�ľ��\�}O�,`^�����C�~���B^����粯�h�<�/�"ѡ��Cq$�Gu;�u��aH�C�g��˚E�Мɥ9B�W��$�&z{G줣<�L8gVo|xGa۱��$#U_��hX<� ��>+N�B�lZ
W��ߎw8�cXx�m_�Nf�M�Om�PT�R6�Kh�VdE$�6�Dӻ1��್ؿs�j�Vy���&��M0�n�@\�X�b5G�
c| �<�?y��0�,����s7v�?Ԃs�v����?��_�O�ד���Q,	��Q;�W��_��8Y �i�6�W�b��7Ꙥg[s�9lE��{��mtC:�=���wJK�h_��+�ێr<O�0�W�uۇW�z���)B��&DӰ�tJT+����k-�T6��v�z�Զ��0���T��{��C��3��G�����w&ڢ��;'�0��<l�>T��ŀ�'?a�e!R��@C;׍WB7Cz���EI�ѭ;8M��ȶ��f��ƑU�>[�S��C��7$jB�	�]Νe�\��s�s�0b��F1����U�!�IV���q�VU��\�؇`�.и��,�c�c~_�%����<������eͫ�a~SP o�y�QV��B����?ЅG���_�j���V��"�(Kͷ�&~�1_��k�*�9��Eyn�\G�+)�gtn�+�\�@��%�RQL�u�}�gű"���Wy՞]	�yTN��#�هr��Q}+q�����|򥷋r+`83$#j|�8׫?�����b�Y	�L᝖+x��v�e8�#��d
t����"dZ�Iy��K�~����,�/�dQ���Y⧈��W�����S P�6����n��b�%f����|��i�#),��i�v���.��p��M����â]�	u%�^����~㌺u)j��$Vkd�r�wڜ�i=2�t�B�{M���4���i��A����0lտ1c���
g�8�$�gYm� �#�/q�)򥦅I����+lw/h����b_�g�قjP����{1�v��x�� =H���&6<�,|��4X��� LFԘS��+����8�"(�:>WL>L�f�3�2���ɶ�B(v���D8�U��N6-ޢ`���Ϧg8;�Z�����𴓇;��1�z�F��0���r�ԗ�Hf>��񏜫5;S*�mT�R�(C5�YP(W�SfA9�R�}B�������2���+���xk�J!f|#o���������{�7&�EQ�wl.	h<�r,Qa�R0GB1\�L��(|uh���B��������j^����$:��Ƌ���mz�E�Y��)�#.>=�t��b*d.�l�e�hJ�:Xd�����j�jT�W����2�O�W�l�a�%1�_PܧFRZY�;H�����8��qFV�MKi^1#���%�&� [� ��?��,s4<�Ca���o�~����⾩��$
Hs��$��@󊍺��U��w|긑�̚�V�O�a�H�S
�J��`��;%V�L��!�g�"��Yt�Ophqб(:	���'Q¡��Lq���U��(M�N̓a�uu��+�:D�@��!-�:+�s� y�5,?}=�B��i*m:�����z���Fb,М���i�NTg�J������:�]`��H;�%R=��
�Z9kAwW�� �1�)/ͩ�-F ���&G7�](}.�r�?Yރ@��9�N���C;)�Ӝ��3�0����?�Pz����qN��6��a!��<}�����g��^���I���|�RA�p:� z�m�8[u^��,	ف�[���)�Peh� M��s�b
�<d��/F���n��_��r����$�@JX�2���^&XC~-:�dxe��!!��|��'g��r��}
���߮ #Ȋ-Y�}k@%��M�E��޺�v�Q��HBM��`�5<��A��}ݗ�E�LH������*TXB�U�xw�'hTI���=q�>m�K8�{C��I�wIV8��bϗ�6���XB��9��Zu��'� ��V6v�: č�I&:��]�_q��'�j&���XR���0��X��|�;/q�GLoFzL��x��{:w�
hf��@p�l�V�Dq9��\��ap�!�	��b�oyZ-�'��-ԍ�-jo���h�� ֵTH����ַ�vB�2�y�8�#�+[>Z�P�~����`�fa�! o�)^	�L�}(���F�p����.K��$��.q4Aכ8�B^Z>�?��X��co���ߩP����/���u�dQ�yS�i�qxmz��	o��ru����/�^�����Im�7>��N��������!|C�5�'��X)�)��)�Ց;��0	�1�����Q��ߛ�������Sbڨ��V�h����5b�����W�(]�|�d<O����PCr��K\��jl�q3$�C�Vۦ�W��h��?�G�'o��гq������l�0l�UYUX�k��Y̌���HO����A�*.��Ӱ�������B`�����JAR]�6,m�-ݱ���zإ��E�#��&Ôҧ>^sX���'���i�7���K]&B���h�ҿЯ3�t֎s{�rw"?1�������~��u�<%��]�����tc@_�=�����}@�v����R^�L�B�V� Z#��1t�'���Ay�t���L����*K�R*}���di�(?��lp���lޙr�I�����,2S{�\9����Q?��g���xh�=���9��S��:M��B�ᤔeq��[���rC���}c�w	hw[r�j�up��j��~�E���2m�w���&`��&��C�7�
Ղ��������t)�+�� �cߓ��,2�w�׮c��B]���L�O�6��p6���Q���P,rT
��;ij����5ǌ�V!����%I�_����&����H�:Tm ����(�����yj����#ґ�$����Q�'�l�$�<O�Ij׼�3VZWl �p�_V�}��s���	�Z��[�mp��˂Wo���ͤZm���~�B��C�n�S-}�s�)�y�@����;����]�*�vś�$EwO�.�-��)��V��Y)W%Ā���0eWE\}�L�m�`�>���K� ���Mbb���bl/��;�EjĆ' G I&�^{��Ú����H��!f,����B���h�#��o�������z� ?6���fv�\Z�^�{�6۔����TL��o1q����2CTI�&o�̕�4:N��fE5�մ���0{[���sС�:�hc5�l�
����5>D�w����~f��X�<򷒺��bP}q���,��,[�Z7�g)��@S��iF2���E�ee"�Mh��%���
3hI]!��=W��l(��EdnΌѺ��!�1(�<}��Z��Ύ�vM������7�F�}_3 ��y�4X������x9Y�e�s!p�y�~t�'8Xfk�؞������������_3���G�ջ�T>�\��Kh�-�C�eZ�y�?$
W�����tk�l��L����8�T���`���̒��݋�Mg��ժ{|�I�6Ύ��:��6�_�ya�^��,���>
�t�<���T_6���Pvū+��t�H\
���~2rj�����ka<�6 ��i���@Vƭ�	K�ߎ?k\�D�<5�t �oc��
Uq�3�0�)[�?�5� s��zrߙ�&M�P��g� �ܽ�bD�L#��+�w�1&QY���s-�,?�������HJ�"��{L�4��3��8)Ο�0�%*OJ���E�̿��j}�%(J�a{gqL+�1[�xH�A�1>�_�^F�[K��*�N���$���@坝� ��I��P�,Z���*�s�AJ�\٥�I�PԢ��������ZE�;Ѐc&.C�ט��>���0�^d��2��a���ի��
ۡO#�`��Q�kNH0��@4����p-ڡ4���e07�����oO�"�݄����p�%����Ϟ�_�����{Db��2��}C�[��°Uu�$�>ځQTa@�������J��&Y�<��F�F�K��seo�aw���;���E0gl����E�<#�O��x}��V@ϒ�D.�E��֮8����0���Bp��T���J��`�����%{�����ܐ�?����Ntԗ��C��_dj�j<�`�#J�7�O��b>t�F���	q�:�b����>����:��6�&����늭0j4�|��=i��$��y��6/��_��y�E�2����b�r��I��2���Mt�0ءss���i�Y|����虐����F	�G ����ū&׭,'���r���k�5,1�p����
%���tB"�n�Z��:�Oƨ�'5�6
W��X4��G��b��1Z��Q]�th2�(n���%@��9l�8���9��h���/2��N���^��!يT��l�P����]k��ʫKگ��u�c��	x�oo�5mo��Tz`9j��R 6[`��v���#%�o�jՂ�c�c:��S�w���Q	-^����VM'a���wi���|�qߏ���D�"�piO�0w�U �M�D����)�����M �<0�]&�.���䔍��
J�U�-eG&���\�5�`ũ���Jc�z_9&��eWSbO�ڡ��z&٧z��=�V#�q��O+#_��+�x^G��&�=s �6\@���������Iq���q����,	6��(7�/���-C���*q��_L?��i42�eAN��O{�+Rb���8�I�v�.�; �H ��J$��շ}=e��ǩ�p$�.z(F*y��i 3'8JX�����z#�J�G���L�z=&��j<-N�0���"��36Bn�<��.+���]��Rz���;��}�,;���n?&�;�M�����!�I7!YX��x��X��eJ`1�-��@v�ϕ,�
�ܑ�&��W�k?��z�^v{�,+�8�U/��ˊF�]}�K�A�����W�,ԙ��!��%���kFN��B����R0�6rz��}��Ͷ��"a7��U�w����QIH7�F�'��K��|������f�p�Q�|#��v�,/s���	k[9�[�#�_��I�)�9��C�d�A�O̲C������rc�P��ρP�Q*f����mY�b,�n�F�}[�]^F����M�V�KT���Y:��b]Rc��wć�+��a+BRܰ~�X�&�V�r��?��?���W.[.P0Fw��e�r{�SdN���ԛ�ì����zR�A�n@06새M���:K�����/�u�T�4Y Dc�s碣+M�eO���%�yi�\o�j���/�;��Z$��d��4�辵+�����rNU��D�D/"��t?j2Ld����}'��"B� 8=�b�˨�����������]�I�`]���a΄ �����D��k�t'h���r�WB霛��>�;�п�B�$��hd�|��ƴtņ�D�������ϧإ\��D"܍���;�޽��'�Ki6D#�ί˿'>42_0ֳ(�k}Zt�(^p�n��X���;�������툡�+�zD̚<�X[�qKL;S��΁�In����Y�':1f9��%2�4���*Q�+�����)r�ؚD4J�+\d� ��E���3x4��9�%�jӳ�4E3�P���e�_y�����'� �[۝>��ݿ^d0t�4+#�ިX�ANs��9��CD����$��<��`�H��1mK<~;���w��U���E�B���	%�:����h�b�=�;*��rY��U��3k�|�R�T����$���r!���q��O���"Hl�Bw�N��c~�L,8�b�������0|��N�kА�)2�cıB,��,MSsT��� ���	2��.'"���^�H��h�B`���sn������a�Эֵ���	^)_k��S~.e��XAd*g�5	6c��mX�I��h!�;4T�#��G����c-d"Eb��Լ7ۣu8��S�F%Hz�>��TI�R>�w�-o��)I�H��`�-ڝK{aN�ܶ����c�b��᫷Y� 6-�]�n�0��w�m��J���g�Հt�<t�?NV�ؕB��:��uu0�����7���k_����v�tl�;�~�W�NF�s�u�/�z�_���,�YJ��nq�	3}ϊ?���C��?B��F�0��aN�-�C��Y�S�4��Y͇��XX���p����4�c��h7�،�Lʕ*/6�Pl����������Ѣz{���YMe�HW�c�hm����H��ݥ�o��k��o��r�������/.�{�>��@�
aѲTf%*{�1��E�ݙ���j���f4�P�+���L|��0�d�1
����������4]��J�A!�.o��b�J���.x�+<�F�V�9A�g
\S��!"	H4������m�`�iD�h�T5�D�1�K��Gq� �Q�GΤ�dk�:�"W!R��ħ~X?��|��&KD��:�^0�+`�Ϻ��Xb�"hr��2����~��3/����`ؔ�/$݉����. 9d'���s=BJ��zn�HJ�^I�l ��D�t��D�%���0'ӺѢ��|�V�?�TB�]�#� 9�i�ϓ�P�[.%ǣ��� �m�Z�G�=ܝ<��9Tr����=�Xȱ�u�-�3-݁��m���)�e�[�/!:�������Ի�EGzd��������PK�����^䐝i����sr�0P��bh&� �����s�Hy�A��R��:��̒M�>�Q�"�Y��vO��ˁ�(�``gh�ܟ�-;���Խh"��ͩFq��o�~VwC�p�O`\��NdQ�Z݈�?�d'�׺���P�S?~X����z��,�V[a󮹔%Z  Y�H�j��mR"��{�dB^�k���^�\*ہ��a<�o�:jF����/8���C~갦�X�>�g�Uy�ët]C�k7�)-0��L��Uw�T��e���pa���;��Ɉɼ���>�ةq<+�VU3�i;��Tv�:�����G��9Z!��)�$@�ߡ�.;�-�hC�9�I'.m6�g���֍��ì��:�97u5'm��m�����Y�Q����ﶘI��"�uP�=�'?;y�Y���y �:�������y�-�~E�Z��_�j�ε�a���M���rOpl��ذ��hZ�5�/����U�����hL�]�{�9c� �X�N�u�/\�%�V.E9���_����;�%U����zIܑ� |c�Yv�l��$���vM#��?Q�5�Q	�?�ts�x{#SgY��v#�?Ɩ�s9�qKB���$�|�� �jL�ˋ"��l��l�!�����x�P+{%}�?[g�^~z�]E�N�Ȍ9�T�&#s��Q�.�d��~�+��Q2 �̧��P)��P�V�:$L �Z���:��W��GKeMu��7�����Av�_�9
#��2�倯� ����,�C�:�[M 7y�^j�!��θA���� n1c��~�IFy-��<�حH�;�ҁ)�o`��IS2j��H*-P�?����\�h��F��$����$��*A! H�x{��2�H�[�nIM�(ҭ�����3� X:��`/(Z�7��Z��_�(�6�g���P�-��k/^*�:໦X��~
�����~fa&��-)>]�2YA��������!���}��cg5�\I�c�l�n��Q[؂�0�ظ�F�~E��eI~��رP��j�xtdd̜�9����L�hw��,�#������V�/�uV�Yu 7;�Ӏ��oϗ's�ئ4����� ��Ά,*hh�l�U[PfM�v!RB�v[}����n�GW�]���p��-����c�Gn�0�v����#+������OXM���!of/L�V���k�/Y�AU�`^V������O�a����hw�0�V�#o������z�f��"�����������Z�:�z��<-R�I�a��}3��}ҦU�8p�~S��I����$�;BS��A0Rf��L�r���h�"�������D�
��v?X�5e'�*�P��:��ϯ˝����v��UɄ�OP�K����G�8����(���N��A���eVg�aN"m7���O���NJh�3M��V�$(���t����N�$�l5�28In$ۗt2T?�YpqTE?�c�2�ƳBJ]��c�ӓiO�[%;>
@?
}}b��N���V:���s(:�tL��Q�8_P�,J�BNE�f��.|u�z;�/�`�Sz�X+X�K���G�XJ�բ/�`��Ht?��WRd�H��E~�C���d("-	�ӳ� �J}�>�ߘ*�
x0�z�������"l@0]{�+�K7�U�V�;����I]����r�;�́'�'��u�Px�JU�;�����O�PN Ř������#�[�Ҝ���o�__a��#nU�el�zRm�T�c�4���&��)3�!ЙH�Ŕ�$�:�r����'i+v �]�T>���8�ה�y��5�=S݋���Jk�<A��W���<�^����([I,�J&2�S�VLJS�`�+���N��fPf��	�.UMCT6�hZC)0l��Pl�t�K	�X�i��) ��MK�
�^n���������s� ����J��W5b��s�RR�dT�d�q�&�e��7\FU�q��N��P�v���˰�~e�Yۏ5WF@W#ꜳ-��w�Ifzc����g�C鏭uRyt�r�yv��ҭ{q�M��ڋ��h�`b4a����M8e��Y��u	�9��M(��U��:P���b�=#�+� �c
o�v��:���m}�o�`��حJ�}��ұMK�
f�Y�f,'c���c��`e�T���k!�c��^Cg�N��o��!���j���8m���q������d(]k~`Y����'�XvT�������iI~b抧���Tt�m��9��U���KY�7�&\��6wV<q���F�5EO�=o�Y�KܵR�E��C�R�R}
����
ܾx�q�N;�z_Ƞ�C7�2��C˄v���ų���i|sdҿ����("^�O5�3W��\�&����Lq�N�~�v?i���[���X��Az(ژ�(�C�A�.�v�#���k�j����u&k�2�����e���<P�	j��U�'���/q���]�v���
�"�,��i�S����P�z�0����ڦ�<���,�z�#��.T�wy�d�2�5Z��ĵ���� ��/y�?)�s��!��͏����Rީ�"�A f{�fU2T^ݻ��G>} ��܀��Tu�-6���X��Cw!&�iN�G����Q�3�f�(�+,{ �e�`i���
(�g�����8[�K1H8���2º-�l�k���ZUP��Ï ����t��w�_���$�����t+YB4�h	���c_��?��+�x���TL��g.M ��t�v[\!�Ǻ���'�ύZ��cՄ�6�S�~|�^v���7so���w%/���>��.Gv����hWܚp��g1�*3���#�O��ɘ1sSRgoI����7��Mɀi�IJ�L��+��Z���&}4k��x7�x���>���3O2�T)�HQj�y�)q�Ы�Xu�{�t�աq�����X�"���qb�<H���d��L6�� �8?i�7���h���4m��\G������Ǻ;+Wƙ�C$u���S7=`J���2�������t�1��q�YD߹�t}<�_�}�z?X�	m-f @�" ��׎ܳ�.��l�m��"�V ��t�b���G�5�Ɂ�����C�nZx��{��ف�jؤWHIHR���`@&~�Ik�JF�W����.������Df2�-�
�KK�Ir�E��1���dbxP��SN�z���F�v����i���,I��j�s�Ԑf�d�ѕ%�nI����vh�E擿�y��������ǁ|�^��Lͤ�wm��~�����}�}�	+��n�x2�����	�����w7�ݕ�HCY�	�����s
Yz#�^��7�
l�؎G4�@����s�C����rC�Π��"!ٱ-7��=��v��6̖:�^����u�;��TBb�O�L���ȣ�)���X0�Q� �g��kRɠ�
(���%��ԶҴ�U�.�T�-�[���4�wxz�gK����O�߆T���	M��	 4=�g��,V�8��MR�>����~pV���g�-3�R��I�Z7���\2�f�Bv��D�"ǈ\�PZ�H�h8��<23VV���`�����q� ��k�q:a2wڅ�����oT�J�;��83C�G��x�y�؄g�<4�>�P��`ɮ��O������ٕ�Ϭ��ae��҂]��t�f���AQ+���qg�J�'�0�'�0#sQh�ߵ����DC\d(z^��i�>�wЂ���`8 {�K��5	�e���r�gҟ�N����Ǌ�/��� D���3N=T���.�����i��c2�#;�e@�.�_
�X����KTsH|�&��P��^��^�f���5f�{*T���)M�?]l���՜J��z��d�B&��h��t��HP ��v7P_8�#AB�b"|����Hz�c(�K�� �$_�ޝ'�1s�ٻ�Ge��s��3��o�O������q�uj�Bx0��TΘ.hKuu�`�����8�Đ9�uH��lC�5�����л:�yE�[T����bjy�Qa�.5_�,X�"�<��z����4t��#�֝�}4m4"�$�y���f_7o8N*��j�Y,%f��mu�T�l��^Ž�@�{e+�e�i�͔���n��WFKLq����CgV�٥677ݰlǌX�=���w_���k6p�W�����RH�bmԫ}�Ƣ3u
D��Gs��Ո��Ѭu���,��\tR���;��^���\��C� ���t�=&�gU͕�z��2��
����\w�����yগ�(7���C�Z�Yz0�S��;�I,'����1��"\�|QL|m�O���L�.�"�#��FˀE�)��� "��!�����G�E���T{	-�^&��>�%DVGz�/k�^0uU9�I�����&�+a ����q1E�:m����j�t/<�!b=��{1��8Z�����'@��`󟯞�+�itQ��_(2H�kY$�?ބ��h��$���	v�.�Tl>xުb�@�}#ѥGh�:��ҍǖO��u�~�'�� �}-0����2�	��e�j!�;��|7Ć�.�v>�W��=�.�g�4(�m�Kܣa��2<�c�[kD$�z�cg�j��7Lk� J���Yٽ�@��'�+�l�~
���.�����v��%j3	�k�ɑҪ4p�W?���`HN--��	��d2�݊!<����@/��o�ǹ�����)�uҤ�&u���!�0���p�?�ugP���7�,�f�9vD����~�qnʶ�y������nٯ�̆H�v���{n4���;����6�iR�D�����_k�Ҕt%y��l����Z@��n
+ۡ�@;�a���\mRd�h�s֡�F#:�*�����hv_ ��'ky�ꔛ�D�5s���~��^��&�և��?�T�jM��E�}�};r�'��qJ[3m+^�k�ƕ�2��b�!:����z�+���]Δ�����j��$������?Q�B���/>)|l&]�6"z�,�5��$��?�h�Qr0���;ֆ��+�E6�ܜ�a�n�E�N�.��@p �1 -5�{���1��N���>u��Tv"a����57n���Ǎ���EW]�+Ѝ��/���]z��C��A�|"+�����A��$Ay�-��_�p�z?Mk�cp�)��ӓ�0��s�"��h�Y�9��������v1�.��#�x����wz�P^���N��=��Ld6-uT|��{=W!�6pz�����Msc���A(�]��<!حk�j?��Zud�����{�6�1��fV�K��JXTP �&���P �sq��)�����_m� a�AY"n��J��3�� �>���tC��f��x�2SJ?6ĀoPX�f�)�WA=Ts�,����q��Q�i
5q붜�b�૴���SG��-��4�&�.:�Zi(��C�_'n�{c�O��MS�gX�gv2=�&�������1 ��~H�^�S��Pt1F�ާ�-9�0��<��|�����a��RMժU����i�>���>d�ɹ�h��@��)pY<;y�H
ߛeF;G�ͲA{s'/��#����F+��];�o}l G!����f��{l� O�
�~�lv���r3��%m�" rp6p��^6�R��`�w���:�:#n���Pr��}RN�;��놤�O�`���WP�֪���6>2��?Tw��GH��Q>�Ћ�ϐB���2��o�L!���|����'� 0U�i>�}	������aH?��Z���z�����7�aW�C�H}���[H�.������p���^N�lK��]�%���c]�{���@~�Rc�"*�d�/'�߯\d���.,�˗�ӆ�R�9��c	��Ys9��L�cA��b��� 7)o��p=�H{QB��&.9����@�DyMHi1��!��������!�Q�=K��[��@���
u�Q�g�
ڊY��!��I�`������9�:�">������r���f��*�3(1c(̙1����	
�������bY��J����~P���ud�X-����N��?O��]��_��D;Uj<�?�>$2�f���l�5�{4PϺp}�w���\��̢ػ@-(j�f��Z��\n�,���h����ͨs�.���	F+�à��� '3M�T	]��S��l��ŗOn)�pL�����Y`P�:�C4
;LO���)CЮ1���!h�F�w�BL�+�cv\�n�0��(H\���T4f�Js��kyb$�v�S�e�:K��"���١��/��ך�rm����e9��ⴼF�ק�T6�jn �`��i��A(U�Wk��b"n��;�S���$_6����D�O�U��ʕ-sTW��	��N�I��Zی�aa���X�SE�G��^n�F���:�s�����Г�Nc:�N���=�����S;�����ϼ�r�e����=^n�4�8���:�����v�n}���ɮ��@��2^Mϳ9`ht.��+��l�b�"�_���9�~�<���4i<��3IȮ|<�P�F�e�b�iWn���&��x ��;����m�r�l5\�ߖ�����r�GI��3�dKK� 1�x�#�@/�+jbAH9��\�j�4n9�罞:��̈́��Z�4���U�Ăȳ�-�|�����9���"d�5d"�zQ�A��j�γ��$ �xDH������~�Sx���sk[^�q��U��Z�}��b���-^tR�=����J[�4���ҁ���Ԯ� �T �zv���-��~�6�B�n���H8��4a�v��D@��/�Y����«���`A3XQ4l��-��ć�ŹB��w�	���
����m{%����-���^�tZ��]���9�U����~�;^���%��~16֢ ��h�)�,���t�[uV�f����X��zץ�����`��\lbIP����I�iH.�zXSq��/�|x�;��uX��o�4��|�J��_��1X�C3��ar)����8�����tr�*a�����4mw��Z/�&g�Z����\�#C8�:,a�"I�G�Z�]��c����B�:�Ȥ�0٦,�S�O�j�܏d<y$�-ǭL���_�)O�6�����s2�#��ĩ)PK	�@���a#d�=�߮��5���M{�4��xR�,�!�J)s���{-�W�S��̃:<����NI�B�H�Ai�!�"]�D�'��n��
I�&K@9�M$pQ�_�tX���Me���%�7XF�H����w����iY(��;�Z�jx�0���	��z�>��gVM�jX "�cJ�Ed�� ���a�M?MJk>9ȸP��S�G\�G��Δ$�w�9r�V�nX<�r1�Y�di^ʇ���Eu��ܠx�����M��1S.o��F�,�[��0���s�q�=�_0�$��>M�]97�6�$��y���It8�܃��@rS�2��!��5q��HG�j�vUz��(��|��7p�l����*O��YJ[�tܱk�*����1����PC4���_7�/���]��J0rʒ8M��-�mqhz��s��}J���m�a��1��X�0���%"�<fa������#ǀQ�/�(�զZ�����tUl\��ٟ$��lꪒ�^e�@��ɥ�+>�߹���č��؛�0��˺���c�[���/ב���1"�M���6��뢨+w'|s�_ϳ��Z��(_ۦ��N#���-Ŗ�I�;����}��*?{]ط�v�T�'�k��T#v��<��?�3��G��k��X��Ǆ}���#U�;�E[#f�+���r���)�Ê囑`���J��3^ `! lD��İ
��p{b�_���V��]�G:� *L��������=T�s�[,#�/L
2W�hC�̕��UJ)�5RdQ��[?�іA�y�/���y������BަGw��/e���b���j��{8��W���E�*;���6�k2AD�i�>���ٖLq%�3�ǼV����d[�rK����xe�נ���p��J���J��?���
u�U�xx����0(�����ܯ���o�����~���#B�0��@��H��O=6A��~��8F�^��T�/��.W� � �T�'v��S/M~�5.' ��?dS���0�;����ǎ%#$P���{GB���[eT����ݻ�_���	�Uڞ��P���$#\�+`ﱓ�R�`���L%]�����@#���@	�7�ٝ�m���0������Z����-H�Lk��V��)J�c�Ā렘"0�x/�����i������A ��]���Rߨ���ZT�UN*��u�����'L��ɺ^l�aյ,����-"��іu�hC-/�,���a�h5���M)g�q]�N��u���QS��_K��"�y�3^-����F��I�i� B���7wءZe4S���>��ꙙ���=U��4�g���Q�=_Vb�l��W���� �		��{�@�{ٲ��X[�O�%I'0Rq{�?��88�0p��z}�'*,��мp�q�����ÒO��J,�tT�h8j.^6)5�g�1���������#i��������:m-�z������ZF-<5C�e�Y����%N �(Rcۍk<!�P��*8���cjĻ�
߲K*��j$�4�Ӧ���,� ��p;�_@��m�g��Տ����-�C�7`h�Om��K��O�֯TH`[�6���;R�i@	+.#(���?e�q����~�X����r�C�Ҝȿ���'m�+�ьx쫼��3x�B�n��y�t|�+$Jƀ��x*IP��#K6S���z����^�-_� �\C�W��d�>�EW�0��RʱH��7Kk��)�L$~>&H�>�w\�T�ߐ`ݕU.�ad�k����6���N����p������e��$u�X��s�q/��=q�l��Ja�/�b��;>�NZ����B5h��"�y��<���O�Pj
vP����HTu�L��#ϋCr�O��S��rܔ.8�ok]���b���}F����O��.�� GL�M>�pm��gK{��8M�/�ѱ6�܆E�2�&��a�[&���1iS��+�Es&�e2��8���$����\�"��]8#�S$!���u�!�,�S{�;�}ɔ�;f�w�%�H�`��!����:"??�|u"'�5�dq���(P �Z ���=b���}�5N�W�y�� {�>+v�Ծ�+�T�` #��l�t����FO�?���"�@�+�=�x_R�F�&"/~6�b:�m�M����bpS����]��\Yh���y�����Bzw�
���E�.#�Uiw�=��=47| ���  b6�&{yi6�y�Z��z��To6Ua�a0$b�$KO�bV�d[}��[W��R��O2���x����p���vp����Y�)�vFA����38*r�r����Ti�V�0,V��#��;��hGk1.✕�����~�T^os�� ��`�HӥfG�QH2J��L�t��Hu��rsĲ�%���j �!��3F�D�4?���U���{����w��+��6#ҷo�����RL��	*�]�=��K�b����Id�Q>�Y�#���W�����<jr�>u�x��*�K?�B��W�lRJ��]�ap�9<�uͱ8D��ˠ�;zi󗬵Jyſ%�;�3NDQ��;�+���PY�o�%��hԮ5���@��
��A\����� �(I�Z�H����^h��?�jw\��SvÃ.��@�>*Zs�S��{�ѯ[��''���<S�H��g�Kq*2�Q��'CL"��:lK�`k[yh�
�(ϣ�BR]���0��&$ﮮ0(~C'Ep�����8�2�	z�v�o'�]�Y��D������زR�P��]w�R���I�Lm�~���9k�	�a���g' �Q��k�~}�;5��w��=S[{�����)B�4���s
���Y�l��"�`Ϥ�b��j6{�?�K��'��X#9�ۏ�&�W����{�	����Bz������}C�w�Ɉ��z#�POy�/�� �r��� �����q@@z^�}F�y�2us
<@��"�f����}{�י�p.�'�ᄦQ�@\���Ig����ٵ����cKb�!�K*�O��K�ŝ�J������56��u��l��T�(��c���F�IΫ���k_A�J\l]���x�LD[�Lݐ'������!��g`�pp�����]I}��0�λy|�Aq�i�p8� a/��u�by���}V��hG����ھ1~\,�n";����AZM9������]qG	�;�M���θ���4j���$����7�����[B����a+��ܛhF��YQƁ�B�KEt:��=Mfs�o�$w�5
M��,`+��Tb�C�� f{D�W���9�N�iM՚���T��Q��m���[�9�n����EϠ��5���O��Aq��ab\@���AxG��/K�E.:Q��g���3h�k���h�)�&����:�")U8H��ȟ!����}|�{ *7�R�30G�lg�9f��'���cV@�oMB��y�*D�So�-�S+E��=v�F���g�NVh�,4�e��*���M��|�:,�ҝ-�`�^��bR����~�t�^Ѱ��Q{:Q�y�u+�<Zү�1 h�~ĥ���|��x�2�����<�!��3�;��� 	Y
�^�r���Ӄ��ֻ�� ;"Jd���9kk�5���kvtQ�(�p�8aDV�	=�ܞ�
<߃݊�?^��:a������W(�^�* �����;"�,� wL[8`B��B%">V���O�^�5W�	e��B��֫Gg3=�F�,M� 0}f`��oՎp��`�����܅��P��i�2x	̥�P��&�Hw�rFz�o�EF�[�G�� @�]���'�^�A���}��HDf �x�g��>^���RY�!�^�,x�Fi_�=��~SK��g�O9�v����\��pg9ڇ�,z�;�L�h�iM��+�+j�L��V(WX�����	t��o:^z�*ֽ��P��5�A�XvZ{�N��X�Z�7��������� �H6��H�����~�?̏�@G[�G���1)��}�)�� s��:L~#��w,�6�H��~�ý���.���X�b(�6��qgE}&I���V(�gP�@^�Z+�����ge��7�<��'�=�k�k�>�:�ig�s�\�^��%��8JqU��&0.�(A%��zao��y��Y���&Q5"QJy"(@��F� �y���r�}C���0�iGb�JH���ާ��0J�*�Z4M�5�L�zE�������T
vZ%�C�1��ʡ��[�r�L��xn����]�L���q�x��헢���{ ����Q��"���� ��[�mb/-ٞ1vF��J������V��g��^g����|�ʙ��Z[��{��L�a6��E�G�������4�?���G�WN29/�������='a0�;�~��|*�u�,cf9���9|���|�;�dN,���ծX�V�b�����1T\u�sn�P9��h�z��g�� Я@K�w�_
��+�J��B�{ �ѥGE���j@��h@_�'��g�?R v����,7ie�i��?%�W�O��9�DK����B�>�D�0�K%qyY�k��Jˈ>��v�v�n+�j�B�ܐ[2��SVˠ��Y�ϊ��e��*Z:�ճ��.�1U���
v��o5�I�kl;�dSh�?ؒW��z�f�>=��Y3v	������%fQ8|[Ӯ���1��ah3V�x��kψ�ڗ^�$�$4�JH�䎈K�D�ʁ���|�����ۄ-{�."��6������9>��4i����[��PlT)��ҶC'k!�ʻl��� �Q5N�$iѢ�Nz��Z뺾��TJ�qB�f�ĭ��)!�ӈt�(�fV�-�����?U�7���z@}���s)c{P��)�3��7Z�)��a'�b�|Μ��Iݟė�2�ܶ��䑈8d�a�	'o޽��	�cA�pG0�>2M�H\� Ґo���]аu�Q�S(rv֍��N���z��`w�geb���P����ӟN�>��/`��6x�9/��k(��Hf��`!3�O���s�9Y�89g��OćC��=�Z��[�χ�]�(���l~w���F�V2=���l~{�{���j�
��.h=���H0(�;&C
�%�X�	)�� e� ��˲��7L�[��3';�jX{=��i�3�A��zyE�4�r�X?���,m�6�������AX�����6�	W����H�s'��׉'��Zl�Z�uh����'�+�;��"��2At�VJp7��2�}�ձ������t��.!I�#���-�9�p�����B�Cr�
(�I�r�+W�`z�:`rn��Gy�3(/9y�T�~���!��i�1�@+��#�l<sǘ��x ��M�*��%2�A����C#��/��Ӆ�~�l�2'�+������)6"���4@޼�������A;����tVnew��Ǳ��8<3�r�Z��zb0Qߪܪc�����I�7¹x�x�ӊ��oq��d�>��-bU�$_֚�8����֢<�l��7�dI�
>ޚ'W��������tv�y�)�XcHvjnb6&���H�8��t"��@�pq�JB�`��ޤ�ۜ��Ym�n�.,���^�ѫLu3���
�KW�t�������l?A�jN[��c�:;��n=�^І��v/ٗ���.Y�[Y�}LM�YT5Μ̌���u>��\� �HG�}��q?c�
Q"�)��{W5ʬ����:�9����G��r�ye �f�4�l?�ee���-I�6E��
CHqP��1��~���R��y���z�V�ye�wD��@�
��}�M���Â���b�|����7��j�ޔ���
�W��ڍ���
^�B��4p�"��~���_�6�ї��5N!�'������}<�f��h����?G���G����א6eM�$�Aۅt����S��e�Wg�
X!��X���剟Y���ʼ|Gg?ƜNjCak�0��A��Bu�~{"9��:����)\T���kh��>)ȋu4/����J���œ��P���'��٤}}��)�_�Ra}�w��3�C��j������1�Б�x(��m��S��)s�,�+���U)w����-���*������;m�ݦs�g�k�ʇ׶}!A���U��^���T"68A6i����n f����n�_HD<:���5�����S�A��[�!��`��g�3(t�-�"��3�Qf�S�dO�ꪞ�ƹ�D��8�G�`�]b*�j_L��=d��z���3>U��ñ���^����1h3ݾ�#���\1<�����fάA����
Z����Đ���:��k�2Q���x�W�ٰk/ڌ ��
�?�q�~�g����E�<�o��+���H!��:�C۴��<�"<�zU�����E��΁kC�������̬9$�i�M8R��% ���o�	\��n�J�Y�LL�R]*�C�	zh���E�7�bc�`\�����Z�Z"M����lZ�m�%S��nC�Ia�W{xQ�܆�:)��D%&|�5P�w冼P�AJn�(1�*���\�:����F���>P:���&�f�Ax[�|�3̔���^��RԿ��U�'�/#k
'�4֘�{���rhVIֈ�	����OiV�z�M�d��,���qW�/}��,s@�U�Y��Ӟ�@�;��B�TƝB���I�<aHΘ�Cm�dX���͞���Pf_��mİUD�6&D1׼�2w������n'���;f�x����ū��58s��-ڐY�S55�zJ}1J�4�2����N��ؠ\�~~����1�o���O*"g�� �%{\磌q��O�����"m�#��߆嶙�}b����]�An�Ŝ|�l������u� Y�����yѼ�{)����j��B��"i8+��H|��pKD�ixY��fDi���F�=���(tؽ��c�#A���t�(f�ū�<��F�)�i����7�-SsO�1{D?s��Ue�biN�p���ώ6$ڕ��n�y�����lw:�S�ty3�nᩯ�.2�~b��ݩa^�5�����/������"{��l����o��	G%>�74( R[q�S�$��o&k"�M�v;������5��s"����(A��Vβ�� �±<BA�,;�3!���cyC�OIP�v���0���D�7�nJ�d�e����ĺ-�=�Kj[)̒CD��V��x�Ͳ%i�Y˸�����	�݂H��t�GS����5�[��3w9�m }�H<�SϜ��嶷GǤ�P� 4����0��a7��}���y;�M� .��]������öS`xpicW�yȰFf�W>L_-[�/����ٓkgkp�:@n� 9[D�+@��P��bM�(l�wlYn\��B F^4P��'�a��ZࢱiD�.ώ|oW��y
\C�.�3{9�:�?�p��4��Cm� >Q�%��z�8�*�ԅ�N1�=���>+]
���Cj�H����VS�
�J&����X���|��*"!	�A\�8NF��<sG���,��G�G��4��^W+�`���á���*g�z�yJM>��JZ��}�/֜�GZ�\�/<���K��o��dE)���V�oO&2�!�1��A�<�p�@�W��1�M��!`W)k�5��I��_҆)����CT�%�e�B�P6���v�H6E:�������]�aW���(=˿b���L��D�ٰ�·M���DV��O|��Y��Ƶ@j2Lȶ� �ػ���mU�}ۨA��n(�
��A��廏wC2��ֻ�֩.��l
ɫno�^���m)�3��c��y�() ����[}���S:�R�����8i�}��4H
:d����hn�Ψa���|�ͽ�
K_�H�rdB=c0���9AB�%ޭ����� 06@.��Yy��#��T��R�R��00E��T�V�0���#!<hV��v,������  ��h���������:uL�h���{���N:�]6�[͵�m�uyG,bKW��V�!��>�څ�UI��@�7$�����T���'�o�P��j�R*��z�`�'�����I��aՈ���jdpi���4W�~'��өw�S��*5�O��_�l��/I�B#H0ǈe�%��'[o�T����W��k���{n�ycEK^Y�Ez��s:�'!Ҍ>�8�)H�G�r KGS�;B��������"��`�]zqO���o� ÅOl}3�YJw��f��閭���������+����!��8?��?�oV�]T�r��=gc\rc�˩3i3q��1����1�r({Q���,@:�Y��j䞵%��d�gU;_|f\ �e>Ry�����E�;�`��h/r�����:9��2�>J�'��f�A���c($� ��q�F�P;w�M����1?�%���s�G�[\z�u����m�ѼqE����~� �U�>�ev���/�[9��(��)�X���**���	~���vn���6"r�x
�փ��9HQ��Iת�w�����Χ|��XK1���C���u1�Z�ծ�����G�M�)�V5ϗ���V�b)r�9�2��Ta�$)�}�H��K�-#(��c`���3	a�%�Է�<	`�H�67��#	EJp�N"��s��ąJ��� O�*)/�c���6��Ã�@�*�9��H�?���>̯M��׽��I��G��7mFͤ��tz��3�@����fLUs<�3zK\N����3y����X��7/f7��gtY"M��&Z��3���h��1��C�r�U)����{��5.J�_�G 7W�d�ċ-�cyP�.�,�i���I�z��F殁*�"�w���#A���4Ó��%��ɔO)�[�	5δ���J5A�y��p�~&:�z 5�$[��Ƞ�W�+?SM�����Y\�� �yF��`*U� y���'}���-���X_��7���u��8��\â/�n㶽o6_�G��h8�Co���{@)"KK�����
(���I	�*����3����f�4��.����om�Ʌ� �~ �X2#����J� ~���M�廭�S�{Y��J� �׆JY���E��E�1���b~4���3r���9�C>��A����8L|�˙����6W-�s�m��)�{]��J-t�����B��H�p�N��+#�ή���Y�5�zA� ��o�	A�֕m�s4��%��C)n �ҹͤ�������um���@�>U/c�����r�b�B���I���q����o����m�MaR�C�N���w�0
3�S����Xl
�4p��lø:��cDE��\-�\L�>��½����Qh|Ge�'��:��dS�\
b��Z���+���8X�O'�LO�����F���=g������$1��� e,�{� �+�%AL%!RӰn=�v�� H4��,pF��1>U�s���e�6�˹��( Gٝ�nI�Eӵٟ��7��/c���o.I�[4^��
����O��s+[!����s���ɋ����a�� 7�5�w�!ߗ�	K�<Ri&�"�%��!9c�oKw-��Rx�����>�'�o@���%֦ӑ�ʹ�q���[�J����Ix�ymq�Mٮ�ua��8���Z�-[Ն�_/n��!!1�j
�ˇh�x0ɀ}>�����/��B����6j�ip���N�-��PD�&U>�-s��.��o��tʋx�H�!�p+:a,"br����-<a|�Un��j-�̽����T�"����K��~pu�?�`��L�5������.��a�iDA��!��hy�,��L�)�e�l'���t�>���a�h����I;U%��^o�Jx\Q���eL#���sU���#��?Zh� ��V{ �	��!�I�(Tr�G`7�R�+�/�Lv!��9�e� ��&�����w��q�݉�����@���'Y�4@vKS�-lF�<����k��/���c��;��/ ������p,�Ӿ�� ߋ6-�+x��G<�;H�Kq�!�g��z�v`��s���_+���b�|W)X���ϕ����c����}9�G�Z$�V
s�����UC�؍7�	��eK��E�e��!dê��¶�4�cx��>fCք�o���f�9�8�ꂙ�Pp�u��*!D�}�y���:���	�~~Ìd2����Rm��i��Kڡ)�vhz�(RޯZFLD��~|�O5R��~o"t�$�� �������Ү/4#1��58���Q;�������Ě��a�1j5��E�Dn�����i����0�֜����9Z[�v��;�pӈ���?G�[�?��Ɏg�Ӑ�.����};ao���n.���SRKʞۉ�n'c}oӅ�[��(�q~�{X���"<�4q���'��
Y*��o���¿6g%��O:���6mc_�$³�	+bʹ����²��pONh&K�?�9oUK�d%	PK �©O"Њ}m|��E��4��݃���5/6�4&���Pـ`�T�~���v9+g��K�Fx��L1���+���L!k-��U�,8�t0�]jUa�W�;��������a��K��:(������-vN�|��"��=J
b�ɠ��Zmg�;ڰh*�s��q<���WdqG�T�z����R��6̯[lxz�Y�	hz�r�F��=���
A�2�-����M\�v=�5=O�5�1���"Ȕ�h��e(6(F����\ה5[X��pM����p���[�@�<�1&$��D��q���N���yd�d�Ⱦ�_����ӷ^��L���Yg�@�]�<�LF~R2ՕY�<fr��;��=�� ��*
#��*�"�5�B.m�;긚��4���C����}����X	I����΋ht�_;�s֬ŷ���5�'��Q¬���>C���i������<��ŀZ�B�K��B|X$T�w�V�I����pu�1�>��X�E�>:��~�Mi�W,ss��v3� �*̎�����ʽ�G�Eqo0} *I;�[�	`e|8�
�u��B/'�$'T�K>�"�k���vɺ.?���i�K��wȘ4�IY�y0_s�:�8�
��~v��2�ٚFz�a�^�|M(��r�Df(w9��;y|�1q������%w0�\<`ؗJL`O=u�[���<�}���&�|!��摽���%ٸRu���O&���͝��Z� ����~M�!]���s~U�<p�;P��X�`B�r�:��j9�M�#Mƞ�F0���{�I�o��N�<<h����+�}�9�8���wz um�2��v�XB}���7a��pcJ��7l������Yߘ��;�}�1t�wi�r.�((�$?֥#�[�~D�寴L��1���n���qΙ˧�������^�i�]~��ښ���zQp~=ɭ�L�����8���8�����$�]�tO<��������e�֟�^~l���K�1��UغX�;f��Oq\��k �'0@QPb C�bPK7	���`�;��b�|���$�Լ�*�?�������$A=9�PF����C�a���J4���,�M-����g�Q�T�K���n��h������#�5G_�����ݙU;p��U�d�
;�Ꮭ��ky�2pT���Zz.��� ��J����`b>w���}���j��F2o�K1�K����z޴�s(�߅mt�0k�ꔵ4�)�����a����VLd#�-� P�z��7�@kK!�#�˞s��J��x����mzm��ӡx�AB@
3�Q `MV��&��C2�߈_����fTآ��)� �A�TcD<��l���VKE��؅r��4$�����r�-9@Tǝ6����" JeU)ۦ�;Ӆ{ʔ�.SV�Hi���:]���F�!���  t^��pO��]1NI�Sb9���A/(�6n%t�t�u�G(~���ch�mP�&==�����6�^0"���H���1p�`^��w T%򞾫�[�"ZՕ��K,I���1��4=��妪�\3c���Б*M0��s��b6�#�,IL}�Kj<7�j"���I�H%�tn]p�W���5d�⥊����E��Q�L�O���S�V4�X@�W{�efs��/�.�o_<cO������A�w$�ھ����������KE�#�6�|�'.=�|1���)Yໞob��jlX�X�*_��&@FZ��[�z�< �70�"^�@~v1[�)be��(h���#�EJ��;���
Ӧ����+�S�O�2�o/�|�u�t��
�Wr�V0#)��%`X�SF�
[�o���w�o���MET �$�ES%
�|�!�����{��B�����l4G+*����Z qQ�+=}�~��O�7�B=���F�����4w��� )��"�>��~֜[�x�� \�@._p��P[���_:"<\C�<Z�[�,9���;�
XB�-���K�rz��,0��Y�u	�?��h�|���w�`�;a�Ԩ��ڳ��ߒ;Gu{�_k�n�o:Ќ�[1��ݔ%��Ԇꩳ��i+�����Df�ۻ}���2�(wA�n��=~��i���(�EX��Vb�T85�eq��?� ����N�Q<�*���"�a�;nd�aR�PO�Jrr�Gm�>��
\���շf���t?hեm#
!�*��9�R1���b��k�$Q�0�B;��a����xԟ7��"�6�'Ƶ���L�F�ģ�G�%�륽�pi9�qK�E�����|��+�A��C0�Յ������l8��0|����i�|�ͷ����ix�f���6 }dy(�������nP�Pvv1����F��p\��>��G@��J)+T遣U7��Ձ���������	� �Z-��4�4�oT&�{���K���Xd�*���7g,旜�%��g�҅�q��Z#�zw�����>4�$���1��H�Y�l��Ow�..�`S�;(��\���쐃� \<�O��7�X�+����Ly���|��:K� ���t�x�{R;�z��e��L0qob٫"�\����B�ϥ`O2RDg]7պ+��ꏿ��<�*G�hr|X@%�x����/d-�<:%[���#H*���%6��a��7R�o�j!�OJ��hW1�[\e[gN�p�Yꭜ��y���r<_<�YĆ�Z֍�'�'d]��A�S�1���}]6T�� �+IQMQ�<��ɹ��+
7$�ɝ�u���z���t�X8�J�w��r�[��2yr"(\��1��FH�0b��%��������6�K��Ƙ$�2�r�ap�uE�v��އj��ܗ�.r�m�@�mɴ2h��]�ڠ�Թ=�9u��Svjv~oE�!�	]�9]̽wn����R
�e�]+��ŀ7l�Uv��8�!�(V�x�ՕgmӶ �H� �F���	�4u�S��X�,�#���Ow����9T�ڪK DB;��6�ː�d�?�QP:jdM2�F҆��?LC�����]�X����ɩ��(ayI�
>�aT̀гF$~�6�
�'��-�Iҧ�N���7>-r���wK�s�����h#rݥk�x��j[ʺ�j�k�VesO)f��C����Y����^,Mk�i, NsC�I93H��;�m���o���=Ël1��&�o��BDeu��/v��%����?ݱ��yl�у_y�Z6}ƚ�3,K|�������El�Ct�Ė5�����.��٠��,�2D4gh���V%ώ�EE�˜Ǡ��d�?&E��[:i�\*xf��(ܺH����m�R����ڰ��6Li=�_��g���n(�������а�6�E�H��(��,^0oG�����yɫ��腫A,��LR�}��-�6n������������&4�d.�Y�;H������ݜLG����fQ"��v��ϵ�6��U;���e(���i93�XH~P<4�% K[צI��&�@��~wI�Ls�Mrݥ���l;�����3�h>O�js��wW=��-�<��@^���[��3�w�����H���λ�(�"��#�Z�;{K��ָ����Î�x���"ʘj�ѕ���}�� A�%��$�\}�bJ@�_s��0�_�9��gQ�m�+s��/R`��û���G��ԡ!�ti�C��h �d��f��z[����[�G�z?f���
��9��m��ʈ{��3��і��I��Lg�3+CJƘ%�l?d�%����&u�zm��B!A�����*��w� B��+��|N��N���Z�Z�\0�;����Rt\֞���ÿN�UW�`� ���r�]�:���]߯�nx��7��E]��(T96��_��dI�K�[DËh�G�H�iiWL �P�|� �C��CC�y�崎����-ᒏhQ��� g��9����iLIЕ�����0�(�Ǩ󵍠u�6�ΏT� ���U�_�`�Ex�������տ ��W$$1
p?�Qy�����'��Ә{��[�Ү�k���H� �>�p�Zң�E;>�����	����G}�O.m�������1޳T^%���K�+��[�� ��	$�^�5�+�j�i�b��MsŶ��#n!�( �=A��%<߇սc���N�|	L*_7�e7��ٓ���;���L|�o�ȵ����@
����l|���\ft���u�C]w������L��D
���o��� �D�͈�m��ݪ�@����-�B�X�E�˗�Pk}�[F=��n��J�+���y$��B
���N_m,P�2�c��;��,�`�������QF�Az?�-��g�M����&;�~���Q|J(������m��F�F���P&�S^�v�%�������9�F���
i>2}���0A���%���e��gi`�)\��euoҎ~�Gq���rBȏ�p��@�&ؕ�9Ǟ$&d3)�9\X����m�Z��4�3�ܣ[�o��wڜ��s����A�i_���\N��	m�}�
�C@�JN�O-*����u��/�Q|Ƣ��D?�ST`��^�'�{&��R"=��ym�O��k���M^�s�+�m��I.��\�׶u����k�a�샨��G�7�h{	��zR�`+4�R_�Ի�m�3f�l��'���:M�$k�d�#-�%]6ޮ�~�ɯ܂��I6~�###������[}f";�I�����S��x�o[���sCv�R����_��꫹�£�޲�c/���]:�9�#*��"��n�	�>y�������C�7
��q?����{\��'u�4���筢*�/���<��4��ohs����)��/�8�Y%��=�}9[�ò�dh ��FȚ�FAH�q{��Zׂ;Gd�8�i�^s���.1��tIap���$T��~�}4�q	����KwKt�q�d�eA3Z��L�R�A��׍,׺�l�Ǐ��c֫ �L�/_��f�7��`_Ί�,n�'��}ް��i��#��-7�O���,�����iHK���i3����߽��JX�mu�R=D��.U��7����<iQ�3�'��.w���c�c*�7�鴠�B68�&h+u"ãG���'Q�LD��W�F���2�zc�R�[�Gz�qJa��b��|3ބM�gc�h6�I)b�� -�jf+�b�{[�x�T���*�9�����uV&�?i��7|α~<D��m{:7΋��J�iXR�Jfƽ,�Oc��=�����t(�h7V�������p�N�����Ƌ&���d�΁t�q���ϊ�ob�4��Rd���Z�0�l`:[��]��ķ2� ��Lk�����,d({,sBu���E1��~�=������^�U�G�ӄ}�MZ�MXy]�r��S�)�v�W��o|�����>���bx��>Ĝ��b�7v\,�x��O64�Ӭ�,E
R���n97ܑ���p?�}�1�s�-���-��%���+
|i��/	͵Y�b
�����d��n΢��(�̹om�!Yqe.`�^�)
ۿ��1��Ȼ8�E/�e��J�5�Kd��O2B��G�.Y���j�xG��53ҍGBC�ތk��P>
��j쫗���Q�U�~��]*��+��N�����(���:o5�$O4�s���ή��pZ��kɈ�a���k�T�ϓV����ҡ��x�7�qip\��M�V6R#�|&�P:���X�I>�F䃥p 72������~��+EuK�ܢ���Y&R}�GbK#h�B?��[EP��?0�Ƨ:V��(�Yq�)7xq�) ��u��BI�e�d8��� W;�y��+��ƥ�L�~���>S`����͂������}��,(�7f��$)O8�yʍoI��c%�xqX>�����C��7�+�r�;���\�8���>Y�3J��]�>Oe�Jyŉ��"��.�l@M�!ˈ�@�X�Q3�8�$�id	���<��  z�`������
=�qI��I
�'�(Z�b����=Ef��q~W����@i��T�_���w��(�(���cKV�0����s�L�3B)t��v^�'��H�o��,��PB�qCM�Q��C�&]�fX��02j��{ &��+�����h<�4�Գ��`�F%��ҿV�G�
Q6�$7�I��1�c����_.d��v$���燈�E�}���ZA�η��j�֑���n|�Ő5z��쐅��L��ڎ�c�r��!���"^��I	j�P(E���2��R#�荾�-z�̿fe�b�vDX'O'�aKO�=��n)e,�FT+^
v%U��?�C��_������|�_�8��w��p5>��ilډ��1H(ޖ�L��{��n|��`�6<�2�aB�ݷȢA<��0�|(�w�p6�M�5E#�s?:��<F�^ֶ��[~T�y���-L��Y���z�D�o`_�-�I����_C�D��!��gVr�T����|��~�6�cWm/��u���ן|dlY��O����K�����0��$�V��L^�}��G�+�FY^q�8�v���,M���A����<G��@Z��AM2M�v�uJ��d���n�t�o�)�*˩�
ت�+�''�G(1���6P����j�f�%�;�ϝ�K�]<� ��=-`D�KQ�5ݯvn���K�*�^㲨�y�޲�W�c�Cxှ�A�v��SH�"5���Ď?M���5���ɧ3�k~�B��X�.�:�A �<��tk����g��b�����%8�H$�U��^͞Jd&b	��̚׷W�a� '���'�t1�T���~��"��f�ؚ����=�x{�����@E~C�AJ@J��{C�R�ط@iX��~	Q�u˃%6�>_�_U�<��B��\H��4��eg����
B�"W�Yؐ:*L>��Xee�X������"]��Qr�']��-�i[�2q唝��#Ѥ�A-5��b	���YB$S�c��3��#P)+�yV�'.n����*��ѹ��h�8>Ư��}k�?��e�*��r��O���G�8X���l��!H�K���%A�tL��?���*����f[-J���V��t���!Ѷ�TX�Ս���N�҇��`b��0[��笝߉�3��c+�Xށ?HK�͛"���i���j0�-{�(��{�նIH�J����Hi�n���<┴�T�2�d$�DRҦjW�3�#�
ʕG*�'��lܻ�j�&U���:��+��x����@�O3�f�,�2�#�>�� j����^��&.C&�����[7G(����Xr��m� �ʘ��C��g�_��?���D'�Z��;��*,���吜V5cTqn>�r ����U����䭌_���#���/O�HJ5��M�2㕄���L�ˋԌ��F/m:G���\7�ݐ�`��R-lO�vk{dd����F�b̪�h��#VL#��Q�8�b�I�s6���
�>ц����A�;'�(L%�\� ��zՒ`Hk¿�clW��rU�9H�¬�i�Z�;qhoɁ�ש����(Rm%(Mҡ��_��ٖ�Zs&�*�-xp�������=��x�=��;�!�T�x�^�E/9sUS��gz*w��h����9�
3��2�[�H	!����׹oM�r��~}(��;(P�˿�VF�iȝXo�3��jl�£o��	B8/�od����:�]W����m��Hi�V�=�$�3��tn1����R,�r?����KV<in;�<���.�^�;�F�Gt�v�&��E Zl�7���I�n�������e�&le��9{�|�L�*���~����԰�>��饰l������W>�or����J	�W��:�	���sDO&Oo@B6�#2��4_ -���[�
��evw��=������JV�9_��J�B���r��+����ne���P+�xj�^=�Mj?Ѳ����������=dNL�e��=���D��"y���H�`L�V	���9j�R7���$ ����L��WG_����{�x�ޭ���]+��o%�+��՗J��v㢋p��rm�S�9���tzn�֥Ze���ʳ֫�}f�ڽ�z��1�~��'�N���xs�PJ�u�.ٛ���U��ٴK����o龵4�}�cĦ�'�?w���y�k�P�hLpQ"�ے*�Q��<��LM��B��,�F����������N�+0��h����O(~�:����Č p&V2��b*�D��#;���&�k�#@�>ESd ��	���~��T��90�x���W���q�K@����c.�@d�jm&[�L���Җ+2n��Ĳ����f@�C�������L���{�)�����9!�>�4����o��Ǹ�N�)�9*N����s��)Q�Ȏ6F��,������L)��o��16M�^���}�Mm�Q���5gÎ`r'�i��i\�g�B����I��X}�Ĝv͢�w��jŰqzǊOf��� �2F��X�=�{�>ԙ}T�YN��| �������@سW������m]A,
Zu��1��q '���;��]Rlj/�	?wX?w��ql#1����}|]<�I`�8�������	���EIF2��"?�_U6����"���*���4��B�����V�e��z������7�[�0 ��PK���_w
��t�֋n���q2u�ѕ����A�x�S12��9%+���d%s0�K��nu�t�m{n	���+�9�D\@Q�Y��;�%�G�fv���5�0��A���v_ 
�g�hQa�p��.��2}���:�,/��{[79��v�q�P��5	'۱O��o�hJ�� ��R�s��;0(�X����g����b:{;!���{>櫾V�S������A��)y#�8��1�T��&�J��P(7~6NV$\���Մ(���֏���m����[:��!���X��
|1o�+ҽ�Z�|�Z�m��_���#A^�$�X?�ua���-|�=����)�k���g6��+�jY}�}�ᖀ���@6�7KL����tT��sM����˙�0���yR����Pяp׆�0-a��H��k�!u\z�r��4���5	�1�q�{3l��W�朇HJ��:i�H��	$l��I�A�Z���`�o���g�-�BW����N��s��VWH��T��6	a)j<	�cL�cw}7BJssF#�2�Λ�q�M0�ۤ�R���p�L/�׷3c$6������w럢x�}�%+oI
敜zs��L�+�����Ѷ��xVqtaP|��F��&�
�]7#J�׵ɼbPI�Kc���롪�*$~^�,�k4e��A {�� �� F�~S���.���������T�,��o�lUo�h�O�8x�AJe�>��
�F�+Ó�:h�TG���<�qJ|��')N�`T���x΢D���Lmn
�ub|��.�P���Gj�^�T��lu�IgS��pN�2N%������!N�>7�od�铕��%ɍ�*B%���.����nx2�{w�ݶ���Vq;�H�=:o��۝ ��<��Є��v��S�⅕�ʖ��_����{�إ7Z��S�QT�y��i.�r���{l������k����,aK�w�0�x�	�P��yAjK`��2�H�mq�:}I��pn�逨�ǧ��*PV��A[��b����~�Ѯya '^�3��{ų�u�R/O"�ď)��^�ub�� .�0u�\qUg�� �6�.s۰�I�"�� ��*��!B�1F���|��
����Mg%����HM_�	'%��k����6�OW_$A����d��Z4���؜+Q�Y_�?�����r<+�og��y��n@���	dͨ�,C�Ӎ+S�ϖEQ�s��&c6�
���a�SXy�&-l��F&35骱:m��~��~�~y
A�F��oFm%w��JJ&�w Ȥ"����޷�"Q r���K���#��D��R���eV�����`�
'1�`a�T��S���ơ������t�Ļ��}|�%v߫eX���NH��#���_�3t��)�(�R�n$:n9���Y#B�y�i9��s��<�
t:�I��΀*��0�O�l��Va.����09GENd�~ �UN-�t����r2U�2�ç�Ʌ�p��S�.��R���ك��:���`i��֬dh��f��\ ����m$�J��X`$�x�=�Oy��P�jOcg�c�4��c�N���T�("O����[�����r^��XﳡUI�?��F{52a���QO��� d�b`^]~o���j�Lf�]��єL��(6&��jh�m��{*@h�tՒ�$.{�H�/�lQ�(S��w�lܔ��'80ou_����8�d+�hU�,1�X�zk���Y?��%zħ����{EsЍ궶2*�����"^p:Nʟ�t�����\|-�H�X��DWK�u��+��jC�4�F�K�gLĠޒ�Lt�/��Z�94_�������6��mr?����I�e��vu9�saU�%c���@grhB�:3v�T_�,�W�zq�-�S��P!��Vd�,���br�n!�S��S�Y���*i����}����l�fC]�
rz���������^�c��"	�_�`��!�:�U�����9ӵr��G��B�ޡ
�%r��4c��A��׵�S����i��MeT�ETΈÉ[w�K^��#����h�JT��@����i%�?AްU�Y�#�˽�	̮Tm��Om���@_�t����!3E�۫�(�����n���5A�"o�N��������&+9>���" l��5%�	[�����"ߤ����h��R<L3�+at��05�#4���r�g��Qx�AP(-6���[x+��H�^�P�)�B�5�Qц���,�:����.ʵW����s,�`�N�5����3AzWI��wP���z�[/��q;o�zB0��'#*["�;�[�}���t�Y׏y����i�^d=���̰J�	�L3���7���ڂ�)�K�T{~o�l:λ:췻xB�,�a��~�PT@�i���k)�ᧃ�4aQ��_�ﺓh*�Dr�;��2�J�*T�Q30�4ԟ�t=��4���F�ہ�B�&��?�P�Js%�u��	qs�A��n )D��X~0ǒ�b�&���|���(##�Կ{�jALu�=�͕é�:�J1֗gIE<�����L.��V�C��������4i�$6S9\w91]4**��m'��M�|�yo��<���3�9�ig+��B��`-���p��=Xq����G�Y/Q0=	y�1����=�2Rk)]�Aw����T��ZH380��ɯ�%^|(���2:�7��э�g�ӫ��riR?�(��h^WT��z����1��1��p��d?<��3�^�`馘���􁌂��"Y�G=9q4�[\9f|B�Hr� ݤCC\4�f�C��M�[�Σ2��桶�)��=�v�G�'��%�X��V��k��TxC�_�'Rj���y	�QK���Z���9�k�x �;��*U�w����S{�j�=�#�j[I���Z��+��a0�)�4�nM0pO�R��lK�L朥����;f}�X���2���_�ƚ�O�4d�f�lw�yͶ+������l�Id\�>S��4��ځ�0����j�G����Xi�뫯n����%���D8�$��b�ZB��a}ZW'�;���x��ם����H�O3����{G�vT�MC����Iި�q�§5e������X��ۡ}�Ը6�H@.�%�h���(	*������O�F��Ƃ�ý��/pZ��Nݨ� vf4N���A�/'��?/*�
�7�����Hq���~�o�����C|)�a����X�=��6"�P	X��.k9��hОn.U#��l1�O��� 8KtȆ�G��4���I��|�R�GB}=�x.�I�;I��H�13� ��� �lZ��B��c=n�hx���PsyE_��'w�R��
���<	.X��x�6J��'��YwO��	��	q�{Ŋ`N��Ge���[t_�������'n�g�vy�^0üL�"~E��P<pbƀ�7o/H��f��>x[کS�^�)RvQ4C'��=Pkm�*�D4��>���YI�J�	�ؤ��r(`	 ���P�*���M����1h�	�D.}����1�@9�[�ݡ{�� )$a�_��0���;�ԡ��	�A�$/�U92��h�"wS���n��-��V�591��su2����L���Ո\u�����)���ŉ��**yR��� صiC��(����{:n�>;�i-u;���#.>P���<,�n�0��z58Ƀ#."���Qn%�Q���m`���_���R)����ˣ}��@0��l~ŉ���S��=�no�'�w���-��UO�.p, ��}��W꓁f�}���A�ӟz�F+ω���� |���q����T��m�� �v3\��N�W�W�/�7�*,��1_�D�O� k���	��B.�댐���Xc(݉B��{7f�Os<�G#*%��1�6F6�)��	�w=uu�H���=v6Z�ݮ?̽��V|���"�v��p���O�n�����JB��~�k�GJiq�X������󹢷1yOm�L�Dֿ
"E;pp���"%��9��Ҁ��9o}x@�pӌ����eXE;E1�T��O~�(�|>���g"zl=r��d�ߺqM����E���4 �s&�0����]����o�	q�(� �	��ڏ�֯^�m�+Ozpd<х�.�=o����a�_��ܡ���_rۍ��uy��ni�ǁ}���~H���`�5j'$��$HDLQE{��@BrF|~�/��K|�t$����Wt!�v)�K�#ȖU���Ԥ�\ܯ�dU�~=LJO�ϢN�8\L7��"R/JQ�Ob/%d�u�_����ݗT��g;>ܛ61[fѭ]��x��{"v�зR��T��7�>`��b#/)�`"��Uxv���$(��j���
b�i%=-C���F�PN��b��%��.c�ş�g/0z���3��Z���C2��]��1�g.	 �	���_��c:dX�V��5?h�I'Sr*�&���K*���A'@���%�9�ԍ��2xh��<���ց�J/�x��dGqV�t�^�ac���[�:V� �#oq=�������!%O)��,�)���j��H��lfs��ͻ�v�ֈ�_�1I������z��FC԰ӵG�<�Ǚ,N��!���=�7T���_տ�7I6����Ǫ�N��-Fq[����C���R����4����R{፬�=8k������y"���8(�e�U�h�g����	)���$=����`,��c�83����'��=c�++��®�FI<�+&�Uo����iN�ߥΒ]H�e3�Đ%`H�<�;9�:l1ȟ�[������(���ӊ��|� ?��X�B��$���Id��a��������'��l�VE_z���ڀ�3��.RnEp����!ptg�1%�S*'+!lҭ6�>���M2�K9�;�3����n9ځ�~�
��v��P��W�X���$�Ҕ�5%	�v2��Q�u?I�s�� ��`�<}���*f��?�<�I�pO&�DK�]Ȏ�ڕ�)5�٨L[V~��w�Ft�+dnH�z+l�E��fԡun�>�hZ�/'�@	Av\&I�˾��[,�a�ǳ��g�G!E�f,�Zg
�(�o�$��/�����P�%��ܠ����M}A��P8���ӻ�$�(�d��SHv��Bbە�D5/��Y���ɡO�G��W_vm:b¹�x]�S���Z��a�j������?����B�^lZ\�q�\��p���C�c�\�u�sN��uSO~�͐�K��l�k�b#d�}��Q�*�`����Dl��m9��!�9F�2��d3���yI���i@+6"e�I�ۮ�;�3�d(+��{�z��)bI�iM(��t���p<���!u���1���Ŋt��+Q㮥2N?yoaQAK�M��D��o�]�	����U���UZ9:��YFGl]�^<�K_Z��#�������,�i_��[\����a�qTLnF6��oʈgd�%��w��H��u�C�y�g�+}��@֜<�L�N��VJh4�4�J`��y�n{��L1k�m���"�T!��Lѧ���g���Y�T�%|��*g�]�^�������N%�ب�݌7:�;��?*0�@M���@Ac�9(�\�!�?9�_�����Cѝł�����3�j��͋�����7*�Q��Z�o���2�D�=i�sT��΅y<?����_2���։��&hQ���Z�l�A@q��W=��S�&^���4 Rޏ��'�L���4R��^:�n0�G�!n�
�E���N `d������WӨ�o8"�g�K�1�yell�r|k�Y�&=p�ϭ�/h窢�h���g�m��ο��]���!���0is��m3jÏ|t6�zP�g	�-e�轐��	�i�^�|*��@��g�m)��X郐h52D�eP"=ׯ�8��!����ۀ�\�vh�C%�7�ۅH*��A#	��?��Kz���?��iW�Δ�0�����d��a��_��,bV�U��7c�/���{,��FƩN��@D�B8�tߥ={5��>W����/� �O걱�糼rǨ&��e���u�L���1��6���wP��Ou-8PYe8\*�t�Ԫ���~q�t�:<|�V���;ۍ9*�?rg��@z��/SQ˚��[,K�� ��EF��/jo�u?V|�CߞVoe�H�������!���"n��l�j��m�Lڄڑ����FcW���*Y����"��]���z4[��'��6	���r8����t"�y�G��(�(v��Lo���
A�`��ʜ�-��q�?za:�>% ��ߑ˙���*�I����%g+rd|�鶕j���{�A�^o��{��l��f�G�%���I߻:����8}�
/ȣ�r�E(=�B��Ң����Y)I��Ф�
������}ca�����gK��O��Fy ���mᘊ�����
U�U�q#�߯�XcP�1�������!���C�G"���9a�����_g���w2�|-vLa����.�F�w�Z�������`(�$���s[��n_�d�r^��x<��Y�s�s6��ل�wl�B�KR�'v���o)T��wk9|*�2�Lj� 4ɉ�����~ּ/����b�^��������Z�&��ŉG���ї� ��ȓ2WA��OcV}vK����X�.�ZCe�ў�)�"����~$����}�t��d��`$�``��TP��Xj�����/\�,���=�#UMR�x-;9Ui��+��SLNr���
�UiO���u ��"5�B�WHF4�mF���'d
��%{l��C`�3��W�����.�u�
�\�/o�f�����,�RM��|H3�.�xɍ�̱�U���+�uS�_������*Y��(q�j(�6�� �?�Z3�m�J��a���uz��8;e��iP�U�4J�����7f�41b�+j�ɧ����n��
&����D��R�:8v�S>��n�}p�z��7Quf>��	xk=����lf�'y�Ns�Ӻ��	\u�u-���\��7�J-`8k�p	��(����-�#m��8�Fـ�>N�ݭ�]�78�r_m��"��P���SRj�7�����Ulz�&j k�9��Ox;�� %�P#�=s4_$:�j2�M�5W0�C�� !ݟh��/�����������H�/����-2yq��@=�WD�
n�i����R�+�#�7��_ ��*o��)*�r����l���e���Z�����N��X�D��p�Jm9B6����6Z˜'$�һ!��&^�Ǡ@� м����MkUCQ_��
p�~��MH⬖X'��vF��cԃ�"ی�����>����p��պ�pt�YB�9�V������D �~�w�53����K��FJ�R�M�2�a.!�j�:�#��V?�q�:�"�4���g}xR�h)���e!އ��!�Ϗ���T.�`9�i�!�l���.���ײ.�P�o
�(%i+NSlMꑿ�;}su����[�W� �;���X#Y���)"�\�J� ^:Ϣ@o��)B�֭��܌����(%���*:����V<-���	�������p .��B-�����aV\7Az�j+Տ��㣢V�r��&l� C�a�m&�������ߤ���-�j'��e��C�7T�.s�S2�#�$?ѿ
����a`(tn��${5���í�����d�� ��v�~7WWկT��_F���ۥ�{��k��<p-�V�%7x<���w��`�+^�I�Xj���-�H f�n �jݍn�_��r�B}�9XN���;_���k�8Nw2�z� * ��Sf|6DC5��h���8m����x��&Ϡ0H��<*F�KI7�<ndFe,Mɽʚ��S/��7,�w>)�en�t��kdte�'������:~u��I�\���F��?��r�E>�t�J����O&z����(��_�?�Ʉ��h���Q��ٽK��?���k������`ь���{��n\T�;F��C﷝E�c��?��U,�WI��#���q�+s�\|+v1�w�1&��-䀨�t���A9�^���e^ғm���J����~�u�ZǤ�������=�ytӘ���́�,DS���P}��w:����%�[�fA�������Al_��l%�$%f����j�7��Z�p԰&�ొ����y�q�0u��2I H&D�^ўK������K�e��:���a>�������C�?�֝�~r���v��g�Uvcv��^\3@P��O��:r*�	JV�Kc���x�h
+����-�&?Ŏ�3�-���ɄT+���k�q|z���\�Ys�E��l��Q��Ż�����E��f��
���N���� ��������:��h�8P�
��Ȗ��`�J�!� G��7B@���c���#;�Tھ��A�
��~�.X�P�h�E��El���?���M\c��o��x~`��;������}�n�8xbټ/�w�-nꀶ��穀���1X���O�U~����ՙ9f�H�@��2���\���G� k��(���l����3�)�����m��ӗ���#�ې��i�81f�ߐ'���-F��,[r��r��#A��%mY~F��?�'��3��m�5#D� ��KΤ'�:1n��l+��q�F�*��x��0�$�܅�(��qqwM��Ӆ�Q�'|]�J�)vln\˓�����3D��z��]��d�bXv��p�U*��ƾ����Kc��T/�X��'T�(�u��h}0��
�
��fi��v�-��CX��l�o�1��a`X�e8�e���FG��]���x?�t\�/�u�Pv!���֛�A�!f�f��+�n��H�����|YI�e�C�� ߶.��MWM�	`�Z������6�5���A�[�mX��c!�t�D�1�o�s��x�?R�sx�4�s��<i��0��|�1��)f��dMl�g�}��&]z4�!S���NgM� (��������c�G\Q<��>Y$0m�7d|�Y"z� 'B�t��a��^�G��/�r+�?�$�*3��P���Y�pr��Kڡnr>O�:=�좴-�\lw���^/����MCs��D�+���jX;àVp��u�IzQ�{#��!���������R'RCWF(�i:�A�0�ܹ�%����v���5[�X������zg#����'�<&
��3�cL$R
�iq�?��|o*� p�����L�2��g60�iF	��Ȁ��!�}�fQ� $�ے��B�3Qw�t�sd2�?Y�MD� ��j����5�!�������M)ⳉ�����Ѓ^���=�ѱ��;c�O�dI����e	�͓�ٜ�q��Kn��;fa3>�����o[�G��� ��$�^�����jR�3<$c�#�K:E��b4$�x����͎U���D�uS]��B��g6���/-M#v�6+R��Yqa)a|���YE�"��\��>Y�f圵u���œh�0Ŕ���^g�\�.`��!}���G�l��f���(X�ژ�EY�u7 ����ɰdy��	��P��Y��. ߺ�6B����f���ۭ%њ(� n�����N�a��#��)橋��6w�HUTG��hp~���x��o6Q�uؑ
�\��:����Bw��͂3���1 ՘[;�F�F�:�瑵�\�������LR��$���� ���4��y��y�񌪠�X�@�Æ	�ǵ�+DF�5�m(Z�]��?tG��g���Kb�4�Y<n��H����~�+� O4�J�z���Zv���բ��lVd'��mȨ~�w!~J��j��Ņ�����M�vq�i��S4|l�e��g��E�Fy���X�r��!$�p�R���x��_��GlGY�³E��l�.����Uu�L�@�y�/l�1ⲓ��VW`4�1�ϑ�n�X)��*y���/P_W��O����Ξ����s!��R�Z�.	U|u�ޟ�kW�����!�H���(L=���׊��X҉p�T"Wv�)�絬��쩎;#'��9�c���i
6��nQB�;&F��["&����/8��49Pt7�jj�/��k��_�uɭx�53�Lט�����z嶼�B�C���/����8E�'F�xR!Ep) �Fl?�wI�T���!\�:���,�M�Gð�p�l�-�Dq��b'�9�c ��m��f�X��)���� !Y i�h�jo`�0_
8�O`�W��@�9A��a���n5`�թ"��z���&A1:����<p��6H�6�o�3�R�U
�{MZP���] ��p�OF'Y��?`G�����WTh 8�i�ʚfe�{x?L�d�%����|�_�R�V�l/'�~��O6C�F%F͌ՀU�X!���i�֕�m�n��6ON��6d;�FIz�~���o�?U<���j�PL��2� ٬
��R�䔌E�kႋ��s��C��}���@���;��/7L�ؘ!J1�R*�vSR�Fj�R̃h���sM�Yl�ؐE�T���"c��m�_�4!3/�A�g�Ĺ#��\>�e��8I/S��eJ�\^�%P����1yT���=in'y���Ja�v�������W�+����i}�4��9�Ђ[���"9˥A�}�?�/N��l��џbYL��~(�Om���ƹ���{a�.K�e �ŷ�I���'m*)�8�$�R�,�4K��r�Qݧ-K'��j�� d����u�T���ܡj)g�£�28��N=�f#�e�Br �]���؝�](�7�����1��tcn�b��kn[���6�/lW�X�uG���e#T�N����A�,��y��Q]Ԫ-{�n���Z0����%GG�~�A��O�a��+fK-^4i�@��a3Z�,°���?�_���aMU�o�/�j���4�Nd�m�>�V����9�	��=�8r�?�ÈRH�I��#_]�q��6�]�C(�`�<���~GI���`�<;0�q˦�LSK���@�ଂN$g��iӂ2t�F3����!7��:ӕ
�y8vű�z�[�{g �"܉!�8&�������j>���_�\���@���(6sJ#<Rs7N
}����S���@�cbk�h�&`(�$"���4�Юu���9�u�J����!���.E�1��@Mno��*�Z��dM ������4ܑ���r(��Aһ��L,�!���g>/Fz�{e߶(4�B�P=����]b�2��c3��j�r�f���0�D=ꃍj9����O��%����N�`PV�5�6��d�A��b�ְ��x��B�֖6�uu��(��vϫ{�:���4�,T�}�� �zu��!2��a�d�GWQQ68o���H����=�T��{��.#����mio���lnr��7[]9�VS]����9��żY�����HZ q��`f[ʇq
���̏�|�"�27�%�$���k��������4z��X�~Ii�smY��_h:З��|�a�&
�����A"��uc9 -��}ǒ��m�!�c_	Ȣa���Rha�ٸ`���#��C^ք�6���6�XQJ��z��(� ?�t[Аr7�%����,��`�"��T��h¨q%��-_�������^��yf�	��P@�z�U��A=�/v�j�����!�f����	0=�	dx�4��ބ�]w���^� �&���+�e[���D@U\V��gʙn���%��m�#	yiЫ�p�ԃ�g"V��͐	|:�K��:lW]z�}b�7PY�g�Z�f����y�,�:u��0 v5+�]-Q�<R��u
�BU�P����c����*<�µ�	�_���R*x�f���`���`��M�e�3�~�ϭ	��{Qb�-��8p�yX�����	ד|�j{���։��вj|�$qYZ/ �����ъ|MMfBՙ�X�eb��ͫqa�-�9��%ӝp���,3մ1������^0�X_$��+�}Ƨ��`����Ȗ���c��QB���L����1�HA�E)��D�����BU�>!��\+�"E]����g���3/��lJx�Z%�;��m��w���_���*�(�k�X+B��9wpW^N�	�~
�r�T�1bek�a�w��UNʚ�V?5~����eߓ�x�b��<m���j�߶<WF�)�c�iU�a��0�b�Y:sį��س�i����?��o̐�		!.�ZI'	���l۲�C����z�]�ג�8�Ү���"�)^,&�J95U9�SJ�|�Ш�6��F�qn�zz�-w����ã��X�3a����r1��!��m]i.��nBS���T�7��DU�)B��m��(k�ph�:9�.M���'*)\��5�GH�{��B���	�$�!�* }�,ȋ�t��R���+�I�j�5���
+�ó~��V�9�,�݇)Gӓ��f_�^���`�˴4$�p���ݢ	�o����\����>�]�O�bq�p8ܣ���#`��QŠ'\>8*If�2�߻+:4P�����r�����0�AP:~�[��ן$%[����B�f�����k��� �	rTu��46g�G����}��t�|���k��
��$���FI���^�fA4�rp涃|����*d�Ks_�0^.��������I�^�O:�߹�r~�1!"RW6Ҋ�	�+���{/E�,�u3�����G/�-���2��mY�P�h����@{׭7���|����5v������m��$n�Hn~�L���{y������,}߅�����-{�PJ$h�>?�H��=��K-�A��L��T��F+�HT)ظ|��d�kxs[@�рHS����3|�~y	�y�F����"%e^��SM�ų���E >�5����Oki[���6�ag�H�����D�#-�i�
gI�o:_�P�~9	�����ieD�w) ���RG�����K����!��A}�L?IϽ*b�J��f7��8�����h��|�
5dA9�j*�>mE�)Ϭ~f�؜��6ݺP�G���Z�3�A��H3�/��<� �J�mh�f�n1�=�VV��|k��@v�z
K��đ)��:y�&W+t2Jw:5�=B��βo2��uSr��9��_�ӣ����Y��1+dЯ5_��V0� ��c��M :��Bl��@'.��ʽI&��{=PwTX�ύ���$j��'[ǒ��k�t�b��])�G���[�O����XF:�I�S���$IU=@q�)�K[>��q%�k�M���r��K�u��4K�K�&��:N�YD�͙_�}g�z~����$��x|�k��|���x�w �L4<���3���1��҂�R[*���G\��h���4�� ���-		$&j6\�l�v�h�)p�ہPӽ���%��E�>8~�����C���O�����4o�G|en����ad��Mxo��Jʂ��DuQx*�o��҉mȂ�l5�O|����,�m���]�p�����[��sTݤ��/�N,'�;�����
��@z��d0|�q�.���nC����P�Ќ��;炗Y�._+�%,m�,/ގ��(��U��'@�h�� �:1(���A�ۙ��L�Sۊ�%6��B8mS8�6�C�<|{O�ج?ߑ�a�s�>B$Ǔ�.��P)#��Vv���� ��'�������Ģ�I��ԖtP���Vd���Nl���S����Q�L���0	��T$Pц�=��X����O�ƀ�f�D�K��bt���Q/�!M4j	�`��M!���E(
�fj�|�തݢg�h٢"z��p�`y�_�X����g����$s>�̀B>I7[�
K�ZL�Y�7k��_���/��(ɅTͬ�\ii��(��*N})����RdP^��e�|on�DX=��1L�7�����0y�#£0M8���F��:�
rK{}&j^�(vBFϵ��(A5��7�Uk�8��(V>md�/͙�w�C~{��+�|�5f R��ˍ��[�V����hל�7[�b7}���9��E*�S<%�D{��n8נa��NR�]�V�U�~�ʁ~�%�K�W&��q�h��[��;36V�sNX��M�6]�v��'�N�jRLLs�hR���yb���P�Z�B�X^���bh���7L]׳�Y0�}U"u+�n�	/j���V}������aA��,B�v�����
���R�õ_�]��ǰ��~�G����ݼ�]/�s��cA�L��V�D��C���1�T; �9n��N�᳖C�������)����w8E�c���]^|�H?:L]aF���Kp�2.,�A5���rL���m���3,^���c��t�w=\SE�l1q�"�$Q�ۖG7F(���b�!�-&}N�r���;X�K6���V�?�^ʶؒ9��3@}v�(_������颀`�@MK�5l���;{ �_)�ST|2�>��{-�]�s�S��K���Pz�Z�zY���i0�'�tp*�FL��ʡ�u3A�.�*B�fW��s/���2H�V�z�(y�K���r�W�^����ec�ϝI��@�b��:2�X���B~?����bPT6~d�L>BU7���T����e���]%,�B�:>ۂ�a8�^�&�2�S�����Ϟ��kh�����Z.���Ǩudx�&>�?��{��`���Qw�l��^�\σ��}X����8𙋅��r}#�:1p/��N�{tٵ�xU����D��������w�|�A%C9~GB/�c�N�Y�D�.�S���`I��V��VSCm��$��|���r9B?Nxn_�;Ԕ��5�s4a#���<��^ޝ� (���T\�C ��0~ 6�^(?�Zf�X���� ��U`�'%�=�&��X��#:����ʑDC�6��
	��F���tm�&�����j)ȼ�>3�͸��(<�n��w�~
�fJ4�T�X���
Y�03݂r��Ñ,GV�!7�����x|��-����e4��eλa=����x�T���~%8���#V*6�l���������<-�v�8$,8�@�1uwVNn����U-�\jE�h6R���3F����:����$���.Fi.c($�B~J9c3)��5�^���	�G5D����P��d>�s���*�����d��ǅ}�<��h���N��1m[�~�'ǯ���5���G@?��n����y��e��ޠ]���+Pv�}4�:����"�R��M)fc���kHb��In*�hD��p^������3��9��`�����+LY�lNC4Hѿ��e@}��p^�����?�m{�;�G��AD��qJ+`��MX75vB��h'����M��,}-��W�����I4�����ܓ<T����0̤/X)��j�3G��<1%�c̹�c���a�u
!cof�f���$�O�ѐO �|��p�q���O��� B(@�01[���1��2� x�e�ے:DQ��ǌez�b^;�]��Vwr�`��N{!�����9{-h��B�ձ��?�-1b�:Fl�y*m����x¥�!i�̉h��i%6�}\-6����Z XA�>a[���ҷ�]�r��Sa�Z��ƽ�ʠ�M.�x|2{'{�8��w�9:%��R��z�k���A�p��ݏ(|��Y�\�S ��_*��8����t�v؏�)X� "pM�=���<�����7S�76� 'e+�!��1�\ϱ�g�q��U1���<�_݀�����y�[�9��}yT3 ��Q��`��Vb=��"l� ��I���B=We�#K!�b���f�t7��Ll��O�$
~J���x�����fA��� m _��mkv{*�{����T�\� �����W=3��fI����TWBt��uy�3`:]���ye����0��Ҥ�0o�$�Uއ�|:
���Axsh�8���(U���Y�g�31�>B�h6��ƧP�sMG�>s��ej�>��u��E !z�:/%ݘJx�<Z�_����z���� �>,op
�"����7y����3F����{��>���YC�!54C���@*y��_|�n,F�.�([Q�-:�e�c�u��[�{ ���K���v
�eDiwD��0?|0m�?�������1W0�R��uH�2
��dl1�����ulJ�9"o�D��[�U��g�kf.P��t�6`}{�.��-A��?oG��(&�I�r�(�&�� ��#�������}Gp�ȥ���3����>Hm�\y���X,Z��S��J�I��� 7l��C�+KL)�"~��1xtdp|�O���
��x8�<��wcM� �}݄�:W��ЅY"��k�bNr���RP���Y�����b��Z'�)g�M#3�#��C��L��B�]����Z��8jpҡA���C��?��j'�N�C����ɳd��¬�"Z�f{_:�G�?>x',����5�y	)��Fo9�z'��%-"����p�acAKtet6���d��C���o����(�n� ���Ϻ�n�20q��ؼ�\�R�?����N񋵎��Y&uᶭ��(���}wm��0�jSzx�%��l�Ԙz�G���w���=�dF' ���=�?RU�S�'�g�ظ����+�Cex�:��=�K%O>  � lı�_�V{��"i�<�i?��OO��W�dP`��ĵ�,���n.�Hl�,T�ex&�11���<z����`�P/C
��H~�6xT8�M1 �o��!�NuK�`_����V�@Um����Y���/���ްZ�h�������(���k�ᇧ~J��T�����S��X�tm�8_ɲ�rI��d�����gc���Bj�i�  �pD1��4�Ti�v{��(G�����Dd�1�ŕ����m���hȞ��P�u�Y��M�AM.��ڣ�:b��gL�M�� ����e�z{=ĺ�mv��q8��h�X����#;u"��������-�Z˿V=m�C�0�Z�E૳jW��>��؈`�6��"q{P����k�i�Q���j��{��;-�>�#���\VD'{�vTM�oB�|+��hN��@|����R�ꬳ�{���$^eD�����p�O�z��XZf��i\�� 	?@ �LV�÷�$�ZnvY!x�@ɖ��ʑ��Y���Wy�v���]r J�0�I�.7b����w.�)$4�.�S���J�1��ؚ�sֲw݃1����-��@��jΉ��
�P��y���( ���luD 8S0H�cI$�_�MnDc�+k�V��!&!
\`������ߡ� VYk�, �ø�����NW˼��]�K?D�А�8/�Tb��)��Q���70ͪ��k[`�CV�ع�G�r ���<�"6)�4AvK������Y3FGf!`F>��'�H�U�Z�f֢���QM�x ������,�0���0� �/^|/d9�2���k+>?7��d�6KDwJ�[�FШ`ȭ0�Մ�3�jb�%]	�R�M%y�E��P�j�l]&sJt7V��W�!���a���;�x�N(�\q��2�
����]�v�U<�:�)����q����G3����(�#���Ϳ>�ݿ�2m�_��Ϩ�8�>��4t������j�Drz��b/���T�L�跈��M�EȎ!�J���mį�D�6��W�Df
Q�8k�zm]6��`��eQlz����e�N�Y*Y�kΖц�cU�J���q�N�@�%(>%y�ݫPb_��f�]��c��P-ԭ�+�n�DѴ}e�ѳf�7Qh`w5�����l�$q�ܶ�}�8$�}B�O�ܲ�r�L��)'�_�H�It��:�H��>gd���z)^�\�m�E��$��QR�b�=�e(^WKL&�T#  �.?�!7����|�$+zf$�P�`R��'�iR�rTur�I�n5�,5u ��"��y���Rm,<��'9�n�u3�F%����y�"9�A�U�又O�������k)�	C���^��?���ƨ�Ʊ]�n������3�`��	_V�=��
��(�ퟞ~]X$� �~��P��7bqk\z.Y�7Ӕ����	�6��\���ҟ�>�� q��Hch�O��8H"�U���X�K6����F��`�� ��|>����79�_�=a�����[�3�s�� ]#��������d�Z7�[ק	��?A5l�2l�
̢X��$m�����F����x?Y�@���E���hl(zK���;pA�e0���Єt��{:\i�_�hC�R^+�8'����`8���x�`��ESU� �
	S��c����О�;;��]�����f���2��(�i�]St�vJ�Oa[�,f_��!���������ft�o��SX	B ���cc�00\&>$P/�����%v\L������M���.Vٕɝ$Gb��nZ��2膉�6�A

�۳��0p�ͼ�d�g�N�e<�Ȣ���N�Q+�k� �&�ZŌ�|�:l�_��5| ��j�A�Wb��3�d�b���$ze޽�����GIU����e�3�*����V=΀b�Ik��������|%�7��&�����%�-e,fF� sgu�/P�! ��*s$*ԷXt���~-G��0,��݆}�Jsw�굩^��Q��KJ�	؊��[�s���\n-\�p��cove�L��gȏ�����MaR|���z�\.��賉�D�&��Km��$�a���q�QE0`z2}���*�f����b#���ݬ
[I� OE?Fl4��@L�`��A �i�70O��9g]�����]���������j������*OPDF�6c��I�2�R\WV�i�>���9G�jL�����/���ki���õ�Ls5�ՖC��%���/�uc�8$�pܒ��I���b	�N8���v~�L�#P!�>k�,	��a���������1:��Û@M+W�h���\����]�ӻ|�4�l]o�9�:��>(y7�Եf6,'��=���*X��� ��b��t)9���{��·��`��CW��-=�q_;�ֳ �����_��4i�+~!��#�@��B�k^.�;�ju�0���\�p�J�@�����aƳ*<|���YN����Iԃ�]�ܕ�R�H�Z��W ��D��P����}+]��L�"�Q�$�7D�pa���~�����7~[�"���3p~�߭��v�8�QB
%I�<�����k�nedeJ��EK�?cu����+<y�0��	҈� ��j���9\��O�C����Ƅ����d��:�����?�^��v�=��`FM����qUF�ԇx��Je��e�M箢M�γ���Y��v~!݌O��L�7�0I^s�8a:~��D�_���aEC�4-��i���H6��I3���N�X�]�~�}�=H���2h�{e{�(٫o6�*X�m��˽��Zs�N�!�D�\ꝘUB�%d���7�[�A�>ٷ6T�M�?Z�L!�IF���Oly[������#}Bܾ�1�¥i$)�N{s�5�X��q,bb����̉��%�p�O1�tQPuJ���j���Q��5���u���J�"�7T�Ϙ)�(FQ����I7Q��}���#�>YϮ�J�4��˩��4-6����r\N���Z��{�|���Wm�a#�LV1��֘���[.7�[����]{wŨ�ަd�"m���ZELny�υN3{X$�K���G���J|�U��1���B"�g�v3`p�83SD�:�U�Z�t,(A���p�PH����-�;;�nW
r�̺ꏆ|/I�B��0��Q?�p�4
U8~=�}�|P��O���%S2�|�Re`��T�h��w9�x�0ݵ������Q�L�C��������Y����7�&��NI[�Q�6˜X�P����..=i(UI�<��+d�@<�jQ�
��.�A�f��B;���W5�m�b��	0V��%�V~х8jVϭdp����S�ًw����(?�|�����tTH��n3�����������y䄋��U��������B�G8L�W'O��	�f��+1� ==(� E4(t��L�OX4EQ�Spu�Z�spV��'��r`����aE�7��y�uQ����X!D����B��k�d��.���h?- �a��vE8��z�����X��6�LֵłL��Q6BBC't
��DsK,�~���!N�$L��WBj
#s<�E�G��5��P��o�sJ�����x�<H?����,Q�z
9`�#mB�\k��z��؃����.��·/�\�6:PY�q������RT�,C��ۺ��MF&�-sw���2�/垕f�~ܨ���H���6���k���Et6��	bIs��MJ�,0����2��%C��dBU�ɠ~ ���j���~9�p/?G�O�*=��:]�t����\y]ۥ[�"�mC�
KxR]v)U��61*�X��P��n0FY3�o@�4@�Xd�j�Z.%��S��J�Č��{f!���;�C��PWN����·=N���H���������9��z
�k��1���ބ�Y�0b�0�G��m�ƞZ1� <��xv�p���}��Y���?�՜ܟ���r�|0͋"yX{�"��f�-��(dO��k?���U5��Z�.;�y��N��ɦ�I�|[���n����*m��@�D�6��׮PW)�>�O�� E�i��U��%���-���TIfߒ��&��S�M���e��/�,����J�?�)�S慲6�{�q�dDQ�> e; ݼ˨�)�Oa�z�t,�żd���Ӫ�/'��4�瞐;a��9i&����Q?̘
��'�[wz�����>�̮9�������%�h����|�Amd�t�ҕ6�:�7"=E�4��~8}�HDZQZ#����7O$F��SED/����u�zh>���^��K.k7�)�ǟ�Š��QH����ԣE� נ*Ȏ��v�3kE�yAr��S��v� �s�N	�d�a�)&�:�pɚ��~XX��~��XL�ڗ�y'V�7.u�u��`������د�:�`2������!�i"�i��ྕS/�R_���{p������ �>S�����@f��yLؼ�P�'�(�Q�vƉ�HkD�^' �|�x�
'�G�;�h�N�4ТP�Bo��܆���e���g� P��K} Z���>W���bW|�2֎��p
�~�c���ִK�<:���+=�@���x'�M͛�R��y+o�֯�T�����r��`����"D�vL=�P@v���<������ǋ=���7Iu�4�ǆ��)Bv6F�tq��۳/�A&I�[H>`��iX��M|E�Dt��3�6g m�>ﱍq�֪�y5����e0�
�}b�,�ᩒ-��
I@���4\��t�gڥ��4K2�t��E��vy�;�з����L�]
q�%���hW`]�=����+Ս�~!��E�O>�ռ��[�1�zpK����a��:��T��*cn�����_C7�Ը�� a쀄y��~��'Rc�ca�3����{4Ak�r8Eu����[�2���s7zl51e��ŷ�0+��Bꢏ�g��]�Vz�Ԝf����5=3�
�f4���;�_���r���&i#��HU����^:�/	GD����N��YIPr�о|��N��
!����HzVOa�,�X8��Wt1nC�<�հ��Ic�ll�#E1r4n�"�k�Y(�VE�5 �M�`�����`���8�у�y�f. J�qTq�2���Ճ�FN�$ƺ�av.~��M���^�j� ka�pQi�%MvO&kX�`�ӶBaS����Op]�M�j���)]8��>~�3�OF�T��T�%~��>7��GM�����������x�oup�)��wQ~�'�4�|�& +����}����nd~�FF��-A[�=��H7׶n��%��Q�����B��įŧ��a/��n9wr�L��ܡY���"Uos�������w��~�<Ѯa���\��b+ݹƌ˫�?$�]�bY�����_����I�/��.[�SϽ���NL�{����g%xo�.�\1�'Gb����;�&���g���r?p�k=�n"�����~@��ۦ_-L�Т��/�X�+�Lzg��C�E��/.�b��f���}0���q���9x�P>0�U����#��(�Q�U�m�V����b�<GN��!��Z͊�i�H����k<6�z�����	6���VHB�O6�����,��>{��.����*1���އ]KH��G�����a0�ü����
kfM%�]�>ز~P����寐:��yA�Nʿ��������WĐ(U��'��)�Ɩ��
�
��$�=/�S�������4r۾��5�a~)[�n0)�TPY�.±qa�na��8b{�3%^�oV� 0v��u�t*	�چtE}�}�	%U�����o׿�����?����,2"�Gfc�v�^�b��A��/;����8������Á��˔���ur��VאƪE�skr���׼J���*?<�t;�����`eϒ�jp�r�tN�$���`^O,�g��nl���)���k+I�ӭH��U�G\eI���	ǆ�o��͗4�ۦC��F_~��f=~�x����~p�^���Q�x7�3���2ߵ��Jj�8�ƛ�����g�����h�
Y�ժ'!��qΩ�~�[�">@���Kϫ����o��F���lZ��"��C8�dX� zJ�c��n����Z[�*1����e��03��Kep�{��q��VՀ{
�&K�g�Z>�ޤT�� n�*���&}BQG���?lY��Չ2ԥ뒂��C�x��y�_�u��`��Bya����;�My�P����F���`yrJ�=�`'��: LHX�Q�K�+��wu���k�dx�=�)B`���?-1�R��j�&�U��[�"F�l��+��kƨ�W���	�����6ҏ*n��_3�tJ�=!3��0��sUJ���*'kK7a��� �-�2��L�M��ć�I��Mr��9�5�#l3Q��zrzS�
��C?/����ܟ�;�{���)-��$�Rd[�����QJP}�j��cnLӃ�N�����#�8�ʺ�H6�憧gW�{�Ӂ;��(0��4q�ȧn�3�E�	����惬����.x�'4�C�W��� ׁ�|'g��}��G�C腅���ˀ�G��F�z�e{���|"�������9!*嗋�&�f�'Ơz"qUj�anN�g��w����������V��P���p&��3� ���2R��L#IΆ�vN]�Im֩��	�q2է*C��l�S�>Y�&޳�<�������C����B`�d_���޸�
�q�S�� L�d+�(^�F�¬���C3�w� �����U�lt�pq�W�3���,�'��m�jh�RPQ�2t��j� KLLW��5�}�z� �L�??�b��E��:� �r+�&��;+y&�$w/g.�C<����e*9�-�!�9���� p6.�|��|�IT�3:��m��0�
7t\���ӆ�($��r�L���`D%�j^K�bo���&e����wn�)>5*[ǔ�	_�nW��ij
I�̫�&69%��.u:	*ϭ'4�wZ����_�bc���Zy��5��"�9B�34t���S�oa�^,h��Vt�������Vh#&��wX��F�p�Xsx�P�~C	�F*�%=�@�^N�ЫH!��Y��^�:������H�A=e}eP�Sl��Ǝ+�#o�B����mr���)�9���w�Ҽ���������y@�_+��ˉ>]`� �85h8ME�"!�{����K�E T8�����)+�31�Q�������^�Ɯ!�J�-�o��{5p�>��=5�5�x~�LI����fH������T�H�|DPP��L��������p%�;>˚NȪ��M�h��z����w�����瀀�D,v�G�̘�}�����QX�������?����\$P�P��d�g���J�|U�B!��h;4��J7��<��L��GG�(ٞݯ�g@o�	T����ZR7���v��:���	��R��OO ��h?)�8�3�ݠ!���+Wj����*�?��;��<n���s�}5����g!������_ ��i|��I� y�W���Ⴊ���N���{��C.��.I��er���S~(�g��\�y�9)�E���/����ߝiy𭗨��\�q�xh�	&XJ����ʿ��
#�H.���螬�{һT��Q�U N��e-3�:'���UQxAF86��R��Y��ջ��z�.����Z2��"����XB҄{��tT�ә)�qj�ӌ<���L5��᪍��t\X<B2=1�rm -����Q��O�<�슻2u����l4w��m���24�E_�4S?n�C�*�6��Ĩ� �*�x�/��XelFm½J��c�����[�撸V��D*�ۮ�̛���G�����u:�EP���Ȱ���;���j5�]o�e+�O��������y�|P�Y�VU/4�����ʽ�ɱ讷ި!Gm���hg
s���ЖrNgf)����.�+�.�P�2��́6���sP�MKwj�W�Fg)��/�	J�4�r���G2�']3�ߝgv�^�Ü�*��ǔ�	~��]���耭P�B��P]��`�,��D���X�@����sD!Vj�c��?�śi{1��\��
4���L(ʱl�{�j�5@G�a�*���kOz͐��w��GR�=�o"�O���c��l��f� ZxW�h8՞���Y
����.窗��_-��?��O���C%�L
b���p���7 hA ����_>�?��4$Q��?ه,�v�	ż%ǧ���a�Q�!H�_W}c��M.����.���D�WF�]�P�Z"ر.v��McvF��{��8����~��)Q �i�t���OY�j���ǓO�=:�6tlTˁa���ں�/
[�}\�wXhl�&!����|�M�"j����,pi�]�0����G���7u���e�hbͤ��D|ԍk�B�{����i]��c7LD1�K<�C�'��q��������$n*
$�5,=�P�pqX("��#W�� J��?�e�Lm�Mt��4��c�Y����Bs�6:V4n����l�^���M?��<E��;�BX��/u/��q�O?hGL�����w.�u�&2�tH�{=]���,��z�\Y��b��d��Ϩ����X�ZbGҏ�q|ˢ����P�:?��6���Zf�Q?r��F�*D"h�&�YA3���8�͹@I����#���A�*�X*�y���r�G	�m�/����Ǌ����:u��ł�,N�%N����A ��ԁ�5P; 7���rc����s+��xa��E^�pbq/���3l�Q��FD1.�u����A3��phZ�C��Jŋw�bUVW�|r0�'�N�r�9H����j>�w�k�'����Rϕ�g���V���_��BE�+�>������$xvRwے9��v���#���؅�^ǻ�Z����?���(�r�1��#�ǐEcwy�x�����T^y޺K�~�Y�80D��p�z,D��D0\.�g;���P�KW�-i��U���	������~�!�ȓ8R��R	:�j4?�T~<35B�@_[�/����c]<baX7�?�T�,"�iZ�)Ԭ>	�v:.*��*+кs��]�de�AE�	Tj@ԫ?"�~ο����*x$�ɘ(�س2�����|�[���W�)���(��J��fm��Lgq����\
9>]�=S�)˓4FKO��v2�KW3hE��j�(5�$��Z@�j�zԢ���0p���(� /���Cc/��a˒��!Cn?ߵ⋸y��t�)��)�������b�V�rxV��n�2[���h֥庪�/�h��S3�Q�x��3xq<|����F��Pj>�8��8:^9��;=�f?��-��"�]��d��/@$�k0�a���mi~$9x��)��[�I�X��$�]�iD�[/���B����'��Q�Ih\ �&�_.�x �5~�����|ɍ)��h��ѥ��}ܢ���5���*v�<��p���@���i�Ğ�����Ծ�ٴ��:z���v��5�� �>X!b{�nns�&��JQ��|���'N2^?5�v1����+�;;&�j���k ��ʼAI��Ӌ��T<��h�l�i%�zS�������{#��;�-���-��/���X��^�	[_ω��ˮ��y��@m@"�P�κ�jg;D����E�Qɍ�c��t���{�׮O�&~�A_�g凘��=���L>�=`CѲR!L^;���RI]�4�Rh|y��!V-G�(�VC3��0�F+u{�`����S��Q�P�(��ޝ	��.�	=r�0A�~���1$9&����v�[{�Mc��-�Y�T��,���H>�U{�W���Pw�T����q9�,�.�ґM}H6pNK�֨�h����*ي�u�3w/�n�	ŷ�u*�n��?:�u4ӌ�>S�'����ox$\���Vg/�ֱ�.�O����iP�-)�L��YA�ߡ矤uh�}�Oކ����|�7`��~
E���{�s/r����S�
RV¤�8��!�Q�iX$h����4�j^�!j�Ȏ$x2�_D"�u�ϑ��?l����e��+���SE��J�9���qn%p�2�4em�x���ܾ�)�e5n�L��4�$	�>E�GHW�m�Q�Tक3
�_���V�ի�u����A�b_��--!���op���d�B����B�TX	u(�c��Y�`6��3�����y�2�ؚ*O8}���A.�Xbf�~uc;�65j'��%�v5�=��1n֟����$Cq_}k�d�bZ'"�z��F��ŰA(랙���8!�Q�)n�&�e�O#��{�2jh��D���T����Xk/��t�y�r�ZEV�,S�b9�j�����91�O���G&%!�]SP1��&Xʩ�SC�
�����U7�p�~`E��90�"�p(�,?1�e��Ģ��u7���K[�ߐE����-׈� a��D�Ӣ̥a����rSC�{��n�����_YazAn������6�u�[<���&�g��<0l"��Q��!.����^��R�#�L+�d]����;]:ٝ$i��JiG�]�Z��~H�ҥ��z�h��E�����;2p���{'�����c�p,Yu����(VGz�<,p�\�)�%�ř�c&�;0E�]vռ�EBz95���X��[�p�Ԟ8��V�2���U��������&d��b}�����'<{<���"�諪�s(�m��T�ۃ(�3�+��?�� ��`{Ӹ�#��؆O{Q%I�Xfå%�&׼/��������P����m�%�I�OĹL,H^@ˆ3�O���m��w��.�⸜����}p�!ⰲfd�E�y5/�X۴��GQ�l43�����uD�e��w�ȳ��<�?�r�(���aI���k�6���Bq�/_�6��V��OB�-B��O�D��7-�ɤU4 ��>��ʾ"P�ځqީ���Qx�����[�b��l2LJ�#7Jг@��e�fЎw��aPe�
�_�������`G��� �5�B��θ�f%�
�	[�up����&�O���j��*�"���9�ϟ������b�S�0J��61����q�9]��=�0���@8J:i�PW�n���P#�����l��.�a�k���h�#uL�d夡�+�����zzŧ-b[A:��Q�艴��~f��gm���+��%������#��z�j�H�����5���Е8���O��l_&��Lɇi���;�����
 �l��(朽ڣyE����q*2�~"�X��w���}�/� (3R@o�a�\����Z�e�E� '��޶�,��Zj����J�����Q���{l�/n,=k�u����8�}�A� !�P�`dr'ە	��U���8����G�B6�_`?i�J?"�Z�;��t�~���鏉U��m��2A�̤�,�T�n�����~��Y�i��o-:C\C������[��>�r{����pk�&�x��e0�Q��U �����%J������h�&s�l��M�%����pM�8�.6�ƙ^Y����=[J��`}��=�iE��5���Բ�M��/����'��=.�r3�J�Dm}�(�~��[�ྡྷ6�M�R����V/q�X5�L��6Y4�2,%��n�GJ�=�r�D�(��f�
Y<k����
Ef瞃l蠍73~�;e����l�F�GW�7�ߊ��q�Z���gh����=k#LS�u�AuP���M���"�Ʀ������`!b�q�3)�L$ߕ�cH҈�V�;��m�O-F��V�J0�ȼ[E��vt�| ���Q"�Q(�jѳҎ-r�R9��] h�+�o)LKl��6)A^sS7V%ze��K
����Ԏy����?/���e_�[�}��x���u�aq#����(�D<{���am>94���N�Ƭ.#$G@�Q)V_(P(]���irC�J��"����͕�9n�/�<�^����������O�u�xU����UԔ� ��Kte�peߑ�@�w��a _$��0	܅��=1�����IF��5^t�o❃$�Ju�d�B��K��覜��{c*3�5~��<j?�1�>�͑\��9Q��� !���R��M�(?Y�{�:{é��;uT�M#)#��`	^���v�~걊�����Y�?�^���ޔ�t��.@17{��1�a���\)�%*=��?�j�K@r���#�9 D��+�m�uٿ�?o�U��)���K�@V5����[/|~]3���4��h]�w��	)M1
,9\����c�x�n�u)=�������L�[2!v�uXw��q�;��+}���W�?�9��X`fc�i�����w��r���n�F�4/�- P���yQ����C$�a�a����o<��yr����,�4�70�ٟo�,~�HW�̧ה�b��U���Sӆ�n��a����B�h�T��?��g� .���_\�N⊠]4���>LQ��!�J��:�� ���_K�9�/���:�wt���"~��h#���q�\��9�qE ��[� ��bZ�/U�.e3�i�j������|��S �cq�
���*��-%h8rCW�5��e*�a`��ф�-1�����}F=���������M��Z�d�0��Wi�a�;��m�>-�_�CCէ�L��ι^,���K�A�j�"�a���ة6���7~�x@��#�3���QZ�pK��9�����^{d�C����n7ĳyx���.6���Z�n�y#�)'�Jy�P�(�qF(f�(R��8i�&���g��Q�왆�;��+�^�e����Y��g��\氻�f�� �����c�⿨�`>|2���#���~F�����n#H�9��n�u�U>�3ʅ��ML���Q2�l���l�^�����%x��Q�ܦ��G�Q�%�x4^P�S��4�W��R���1x�3YT��G���Sf���A�A�L�!u�-W_�������4��+��J�	-�	�e&���I�h|羽M�߿�! с
r_��%�M1@��Tf��%��t�������w	�f?�~<��Ɯ�T"�z����v�
W��PQ-�������Vz���a\������ZA�58%>2��w!��tGy�#��肈�L���'ƛ{n��s��TU�dRl�����N+lU
Y?�L�"�~�h_4	m�P9�(�֛;��Q�B��m��<@j���s��NK򤿱���Z�ךw85	,��y�\�5�A��a�w�Zw>�~S�+�t�,W���3�މ�m�VƬ�yԪW���w�R��/���7�(��dI[����u�aS�L��!�(�k�[���qx, �ـד\&�K!�DASK��0&��9��K�wZ�]�}�Ի�Ïԕ���Z��xv������U�ië�����FA�6V>v��<�_?�9)���*�vɳ�z��9�Μ���K�8o���@P:�Ͽ�!ۄ_14ev��<+�1{\���K-C3J[��z��u��jC�����#
��Eq�;)�XV�����������;mpGC�G�˘�M�J�O�rڨ����[�J9�@@�Wy��=�qAV����4D��b@�����Պ:x�%'�Zqq�z8�t������a�$��c��ж�*�M����#�2�F��J��
��A�d{��Q��6Q��o��g����a�-�$o��r���:;. *��9�����x# S�}�ҹ[r���s����:�M��`8�=,0�G�JJ3M��ER�A��z�tq�ʷb�zP3޷� ��r9�Y� цhcZ���ϝD.�찊>�峮�&*�BӦ�N%g�G�����tc�?�3��$�i�	yO�SA�s�V�ãf*�@W��}¡�C�o��x���c�ɣ���8���G]�h�|�\��Dx(4�L��BA�!?��݋"��^��]ӊ�>e�����*��f��X+�MQ�!�2r>�� ]S� N��b��^Ӆ{��p�v��ҙ�P^�&�8�ޥW:�Xx�1�VܜzC�D��#XO��r���Lp%�Tꍑ��.O��r�����cwi:��,�	�W�}��l�Pq�dxJ�(w-�Wa��G�^R����I:�qq�B(��I Q=�F��[$&	_��.+�Coqo�a��mΠ�.���V��|$�9f0_�A�`�5����#�g)qF��^��RJC�'����'fICn�r��_Η;�yAH����gu��G�h�ϠYV<�0h���*�}4�Q���X%+�#ϭ�i�ŝy�d��]��1>FYc�n�2��̳� ��D� x
��,Iqz5�����ʊ�5�����ʊ\�M>����vI�ݟA�
mC��R�S":�L�`�R��@�Ac:x_b� ����x&�s��(����Pz1��t���浶:���%y�S
\��FW��iż��$�D!!�a/.O��s�No� U�N���|�	Jt7+=��R&���L޴��2�������(s�V ��ż�;�1e.;�F��m.Y��>����ߞ,���#�l&&�B2WW�n�� �HP��>�\=vP>�����P�Ȼ5���g�]��`]�!s~\N���i�0d6Hެ6���Y^a
��I��-�uwF��������L��`��S1��]Ti�<O��W+ ���*LǷ����β��L���l��H\���d^���ʹ�l[��tc����Nk�����cd�~�7���_�0��g��^f���ogn"M5o�{��K�G��]����`��6���_�A�R<������I>���	�|e�Oi|���$�,iқ�=0Ǵ�
�6Z�,�Q������S5X�Y��aFk|ҕ*x�'��,x�=+�Ǿ��UL�.�*m������Y�t|���l�p�,S`息�"��xɞ�D4�4����c��M���8��?��<_�yq]��ם��Z��@.O��4{��V譬�Z2�ӻ��9?)���ؑ-CV��Rj��3!�)GEV I���e�$��}���K|"���}�0��8�q]s�p�Ɲdț�jn�)���Vʞ�*��paD���N2���l�W�JR�aq��$>i̒qs�]���Hm=1�>�|'4er)�T��v��z���s"o��1sN���ԛ|X��'���_*O�w�_e2�A�ci�%#���!�t :��=^y��W����3�&��,'(�Q�;���3	�/��7�w$�*B�r�:^�FKE/��ď�uJ�Ӭ{���@�[ni�5�=Ta�����*�ʙ��*x����&2
��$�B�@��Iv���2ט^W�k�]��"N�,"'���@���O�~����z;��#<�w�(4L��}d��2�V�eo�-@�r�N��Rc�i�u}�<p9(ҼtY YB�.mT-c�j%��$��K6R�v����C�8Y��S+���\K0�,ۗ�uԋ�{�-�dS[T~;-��(�*\r����A�M�"(�p-R������BN��F������K�K�:���a����je��Ym[�������,}��ŧ&�����4��`��Ҕz�z/sZ����x���n9s��!��p�2�P��G�_5c?"�We�!�� �7�J2T[k�,C�(u�?��R�Fߢ�">�*Q]G��%�6��b��{��M����ݬZ�1����J�`���D��6uf���_[zoF�W~b8V"D>cR w����E�I��p���I�u�$�EG���t��ֲV���H*��� Sc]A=�_U�@`CS2�>�=��e�5�t>~�������>��$�#9Z�hy�?�7}�p��~s�)Hj`4:��T2��vI�ű�U)��@&[W�C�Q�T~�o��C�|��>`t�<�1�5 ���5�:�����Kl����Gt/��d��N.�KWn��7"S�rQ����FVu$���5B}�XW��#S-�Z��B>.{�����g%�p"j�4�|��6��h�xNO���&�`f���(7�E4��n�z[r�X���%;�#uѽ�4w�yN�/sŭ�r�)��Nt&�I�uv�� Zzb��o�8G��Û�Mdn�:��;ZT��\nb��<���a�z�����?>;7*�H�H�nK����INz/UG�9-,�c���ZOrl�!���{��{Rg�h8�q�4Ld�����lC
�[=����O����]���r�Ӌf��	N�g'�؉7U����>UH?���l�����ã��ui^��?5��$�; �h��x�f��mx@��G:�1���N4r�H_�3�B:>��,N���㳣�_۪@&н����&׃�M��=~NPO���r����2��ݜ�H��:���s���n�Ѳ2����=]�^
��P}��Z�
�������c��m2&���䥁S���"��F3M۴ �:�-��v���7+$u��RS�}���6��<O:������LK�m��I���ooy_��P�;Y�O^���I->)�����R�G�{F!$Ea��a��ЮS��l�^v��:�j���{��1$زf���	��IX����RmsRQ��\Mɲ5��hIe4�8y�\<�r%���>qܾqw�7�v��2 �
>*:^O����~0JI�N�
�&�����0�f�ƃ�_�K<}��&���O�)[��bUfzY����1�����,Gz�j�Ǝm.���Ji�6�Sl=���,:�}wCQ��s��Ti?UA�"rrћ��iwX����RPl�r4@�g�)R�\4��k'�T�WB���PfY��*��T���fcM�&2���fv>�Z�h$�z�6>-��M�N���o��?h�߃���6-w��N��Y�|J�R�QHS_"�GLQ�=�lLz	��OA�Q�Gr;"2��u_	�k��U�\(���x@ a*�c!L~��@Wq<��K�'@sN�f��������p��`�^�v���L�|��(� K�Af�	%��0����6^�7W�B2������S���!��*���}.�v�#��KsX$�"@�Hs��d�lC!��j��h��*��'ۑ;%1�Nz��R���%a���,�ՙ�01��ׂz;��6-������?�@Q��LNs�a|���GKC���?%>�8Ez����p��"}��d��W��}�=p��p{!Xn닐O+I�67!���D�G��������%�L.즻9�ish���o��|fG-�X�s.���,�f5�vp��ΖAl��(�a��R���g���t��D�������Lk�V�^�c
u4#Fy�>��4�.��5�?-�p�h�q��S�F9����;���@c�m�
k澦�K�7�zM�����#V\�t�yԌ�H��e&���e������� d��?s�󢥰}��3a�ψ�D�T�m��!���CL��'�N�9�i��.\^��n=�� ��z�mJÝ����ˣ3�P�S��ԛ�p>�ʊ��@S8�)3V1B a�u&�{��:�a�����Z����@�|�"�9��v��)���3�^���	rP��npGIא��f	[�0���8\d%k'bKӠW
>����H��n>����ɭ3�	LN?1�.�y���렊6��o㪂U�i�;�С}aq�>��Bk���L��� \�4l���*���HN.����C��-e�b�iw������h�+籓`b��e�Ҿ۸ŧUծEg;G_��g���xo�a.�2ޖp�.���z~]K�I:�^�؜Cb�@Se�LLaj\����c�U16@Cw#�GA���e@���'��DH��T"gr8^���Dx ����yv��EL���ƒ�;��|)�SYb��-Bӻ�k��'Մ��R��$&�,nMռ`��N�� e�šL�������1<C�N@�ʂ8 �a͝���L&��)ܴ��$$�'±ٸ'5W1����r�١^
:pB���A�"�.@@R
Q�7�|�/FTO�j÷G*tx��	ՔsMk��#�8�R4u?�K�.���dT5T~������+Z�3��K_����8���J���~5��M�_Ö��o���b�M:�!�$���fB����o�Q����/��2��2��Ct,��� r�y^����#��Q�� �fka%
���H-����"�)��{�<��o7l�������2Z�nb-C`�C�pz�AҾ��fo���?�C$#Vc�A�Nܕf����o��u�����Ke��D\�:>gF� �Nk����E����"��M��-1X�=;8�`f�"{�ɹ0.���xF�g��ݘ������S����
�ڽLk)�^*�c��s2RL/ bPI�o��pd4k�<Qz�C9E�U-�OQz�f� 2���Wx�}&��L�W�y�BΝ���0�J���k6�`^tt=�W?��'\| �Ϫ�r��3�Ty:(���W9A�ǻO���\
�=\̡b���T�F<�{h���\� &5�������&�D0�V�Sק�vW���j�����9H�C\b�Z�Kn��5�z������:=pvw����Y�tÐ�f��`���j�	1����Z�/�[ݤ�У0�6��&�������
9�}gmS�}r��$T&�]G���6���Pe�ã��b�jzؠv�dSL���l��
��0�q?"K1�ŊX���}�ٕ�DV�C� y0I�B듨�H��)�Ъ���/M�Z&��#�(�
��Rq��c�"�tB�1���"@*Ġ9�J�p,�vډ~|�=+�K&6k���=<�yVα0z��!<T&�����n�l=��d髽�̓�R��k��ö0��`���?p�32;���?ʦ�Q���x*�!���W���M�o���V 	=�m���|�JՇ��E�DL�0+��d�*��wʗ���_�*�`���������}�T�Z����k�+����>��_�)x���glU�f t�����/�o}8��:�M�p�����n��t�=����g��Z���E�._�)���i\��Y��X������;�� 얜xE��KX_/P[I�8�����E�(_��g�����h�����]k��1�.f&Q�߭Rf�8�Y�Xnܵ�L�gF�H\����U���d�m,ƆVe}C���ZM�FY��y�dw[��P��0��D<��x�~]e��fEI�{+���j�B �W����,2��`7�jP���2�E:���p���gA���᛿3�����e�SAV��(4�B�N�_L(��	T� W��R��p轵!=V-�)#�R��^D���e��emȩ����~T]�5gaK��}1br���X�<. ��{�_�cuC�{��2���*"˸��H�dt��+PA����ۚ�E�)?е ��+���"��B��q X��7d�H�Y줟ڦ:ĉӪ��B07:H��	,�z�.݃j�-O�R|x��Hu��J �р�e$��hH����wI�T>�:%Y#��RD���8�tʢ�'��k��B��k ':�8�a�o�>_����>������;�Jc��(� ���	��#�e(�E����!gP�/5%՞NN��KH��/�T�/$C��{�{������������H@"�"U+-���T��в�}�����BP�S`�5�s�@�C�̕F��M:;��F���'Z�蹲����[�n�u^�\e�`�'3{�8-�ڃ�jA�=�S��[2�8X�B؞a|�-�};��1iA.�� �7��0��C�?��uB���ֱ	�\��qa\OK���8pa��x�R����b�y���%��T�t�:���K���KzQ�̬�,4T���xI���K��W��R+�������=U��]�I���D�Eb;$�lT���]cW��w���"3���e�\��� �+��!Y�B�4 @�a�8��C�F�|�ӡ�bB�n��22ﷹ�p��ƾ��B8��~	K�d�����\Ǟ�B���5�Zpr�ċ֝�k�'�IO�5T}ܶ~{���"9B��
�c�R�q~�B��)���<U�ը2��Ij�Bc�Vo}枎ͅ2��"r�M�V+�m���{g�@�����5��"*�k�V� �b$�X!3�fFQ0:�����i
&�Q�D�-�ݜ�V�[�t��5��aΜڦG�~���S�o�N@�}�l�P��	5L����Ft��U0)x�󫟋>����a&�t:���*Ly���V�V�������w��"c~5\�`MǱ����̴�f	�-��S�xj�2��@�$�.�9Z�+K����|P�����Eb����B�Q��5�I�U�L�]��`�Sɏ&d�6��� �r-1�e�,�I~�)}�a��M�́V�5W�b���E0V@,�����N���4�Q�rQ�M��i`(�{n�g&��q���zf�"��1şu��nd0p�'���\�YC����������I3���Ia����i�L��g�����Ә������pGH˜���<�e��Ѫ�����U\�S�
?�%�H��L��)_K�dc�/��B
��dk�'�]v/:`�=���[W��؀��<0����ǄML�5���e��d%X�`	���q{Y��V*q�b�[�Kk���M�V|���K;�h!0�B�^0�SG���ti�V�ą�"_��*I�>�������k�W��m%�"Jv����B���O�巠�����#�H�==�b*|=tt%�Q��:��lє��7��3>KCx䘬�k]WUhM��V�^"�>Ƒ@�S�jY%�x߭>8c�z+s3�q��`_Kyo#h��"�`�}}��D4E��;�7<5Ƞ�m�6� ���/H�sWu��]�=�ŷ5�>;)��3�C��%�e�Q�u����e]Uco-Q��I\�1I��A���(/��b��$�r|�=6�3Û%b �k"-a^�ǫ��I���|���ދ��F��|(850����hT�F���E�?���N��	×�
a�L�����9�V���a�b�U�bEӇ���/:�Vy�2���p�.�E{��0��O ��[�W�3-�-R��(��OqKJ�oi\g�N�5U�S{��̭������8q�n�W <��h��0{.�Qm�u�ء��)�~z������5�>.��Ϟ����hj�;k��ڍ�L�ߥub�-��ס��Kn�
�U3d�:�5�mLٌh��l�ܟD��) ��K�� {قʜ٘ƶtf�	���t@ӚZ۫]�:��$���ƀ47}�na[<�5jD�F �>��ӳ%I�2���1`H��h��>bxu�-#��>gs7��b��c�DB�lO��d�
��)��:'C9�2�oG��X�"���į�:<,�j�l58H��,��ք����
u2�>:>�mS��r�Z����F����j?en�	������ڑ�Z���kN���?��}�@)8cR�{˱į?i���R��3ߦ�\�|~�ݡ��c��Ĺ[��Zan�#6�^D��D�FN<��
TA��%n\�Bo'������8៯Y
��O7�wʜ��J�6�x(��v��IT�_xEcW�����C�a� <]�U���D�`vt0R8k�Uڜm�\ZA��R��b!�"�f�HJ�	pM����;�I?�G�%��3�j�B7���	9[�</^�-)ScK�/"6�X��S:��`��cqz�_E(V�4��q%p�v��lLro��n12��le���/Dh���-��v?EǗS�wNe�?u.Tg �#i~~�gn�<U�{P����E��x��Y��`X�	��J�t�p�܋���匡5$����_�3�����ɜ
�줦NV5X��r��e��F'u���u_g��_{�R�5R��th�8<~{��Z����(����*sM�:��<�sn�e��` ���oO�0��	l&%�����dU�!���.b�%ԏL�U�*��q�$�~|���S`��#���x��8C�4�H���K�P
�z.���S���$p�XJ;����DsL�	.��+LL�I?n|Б�(���O�ia�%tx�d��Wb,RX0�b�襎o
�>��Έg�V&���\��S�u��.5��L�E���w���\:&kHq$��'�Q��r��aW�:���)���G�Z�A}��1��.��^B�<
��cj]-O����%@<N\� P�;�o*���L�Qgx��H����	j��rCl<�s�@�Y��dp��>b�~
ۻ��y��k���c��e�)5^hH������̬HC�c�1�c4�-���&!f�u#�0�0N>h���z�8��)���ߎ�L�g2M>?`�	q�Yo0��:�,��Dv�V�9�g�W�� �L�r@����F1ۃ.��*���#�d,���n%6PT�)|�'��H��&�}�	g��\�.�X$	�K7�U��d
���O��p���"?��3�cD2Ƣ��]��/�����^�W�����|�@�:W��-*�esy*�ۮd�$��܊?�w�8>H�.�|��
w���:uU�	���S�k���Ak+�����G�o"�%6��WO�������/���ne~�c��c�ty�gX4��鰬���9gS�r[��ant�v��<)iJ�zA��W�߄��[W1��<�"��hW)�qC�z:8��R��4�y�Mt6!��r�Y�u���ŕ���ʩ�HV��U�����ѷzɱ�ݼ--�.i���W������T��������i@�8��z@��LD��(<�x?��hžɱa��4j��`t%x�I��,ڣ��TYͮ�g�4��n�Z!v�������LZ:��7��?4���FL��.��o����A��D�R�b]���#�	X/���3NV�A������&I���ў胷�;>���R�����X��G��_A��;�TS9�*5m��_:�O�=C��?o�3��J���8��{2���o�����7�/5�k6c>���S×�׆9�Y��hn	ez`E�j��7az��xr'�'��xJ�"͍���!�R8S	�]g�/�0��������4�Ŭ�J���F
PAY�<T�z�$�R��n��_�%�[k�\@wmg���D��ݭ�?�x��
�8,X؎����!㨢\�T�	�;��s�]p'���o<�^+_SK���k�gPho�0��� f�!�TT'lCP����}U7x@�a�SXX�)�`>h���QTDM�qxb,��N���c6�oىr/��/9�M5��aV<B��!o:f �ïz#H�Y�;È��!����� &l8�]����!�LlR�w����S���v]����ӌ=0�`�
��<�X�Ȉ��4q�76�ݑu�
a��'[���w���~{V�s��>����x�;�����+,� u':��47X˺�?~l TvLߥ�Z]N�2�b�W��v�d.�Ѡ��s��3�+b���0P�|���ثk��#|�cO�@��U D���DR�x$�N���škj�'Oه�-űA͔�j������V�J��R��y�޺j��L���b1uxE5�P�ָ!�Q���g�65�.���_ ���;�s)4�r`��ď�N-�[�HK
�x_jS��xH�%�r ���Q|�Y�_����a�y�"n�G�w���Co���j�Pή�ul8�%���Ru��<t�]�Ba=!��yX�I���{��܂�"G�Y�%Ybgѩ�,wp:H���6��'](o�-�B���D�C��ퟰ�N;�N̄ح��ʃ����G`�~:������D���S41�5Z"��0�c��ۊ$�~a�>����Ʌ�oLfat����dD�T\Y��_��	"c�i�A�#`6���J�Q��&Yu`?��C������N���5�D���R�뛒�B��7������A�k���Y�m�S�Ba��ւ����݋4���0��eq���	����i��6�	��ɬz:*�*��`Cd����}���:S�B���@������Dhw�˯J��Ԋ��~�H�MM����E8h��	K%���f�kp�yw.O�{�F����"�Ȕ�&n��@$i�IQ�,��-2� t`��<�tW_�a}��$�p)O�(��Ϧ�/f�ㄡ��/j�k9qE۩�������[��
��t>��b=���1����%���*����E(��ޚN��<��=�cYu���g�9'��Q�ډ��qѥ�a6id~��R����e��J�A �� ��g���9?��=���@ebC+��~� t���͚��\b&��I�ZI�����!A�.>���÷J�;i��� sF��޼�#��W줪j�nvT�F����\W��B�y���:�g�ב����:}�n����dB�<���~R�8���dG�6D׊qLh����ç��M�9���Ned [����?�$�&�7����"�U��@x?ȭ&'��2�*��r�^e/�q0�:hJ(X��{�6I*݁"��E�%����}L�4�/���IR͵��'��bO#"�J�rL�g��+�T�g����+!��]P�jw�C�`��{'M������H����ј��[����ܛ�����O�����uM��j/""K�@���*� kŔ�?$�a<�T�)���%���y�brw��bTHɻ�F�_�17GUo���%����ף�fW�c���_�2�VxE�	�;~8t���7L}Ti��s������ШA���nv2��ʄ1���M@��8i��^Q�7���c��D��`�v�(a
��4MY�߬�:>=�b�hS)��q�����L�L���M^�+��AY$a��ٕ�/�ך?s�`2��!P[	��J)Xy��i�utdX���߸e�3(��\55sǦ�v��
c{|��|q#函�Fa�u��R%K�v�z(V�-'ϙ��)�R�JPA��jE�`�c�2�K�&����N$tv�!n$.��Q�m��Kku1��ˏ��@ &V��A���R���2{��HnR���½�j�������u���5<\]�C)�jr���[?��U_Ώ�t��02]�������_��r���ֻ�u��`���8��P�R*���&�KU	����d #�upG:qq�JۂI���M���:ǵ�d�k(|���Ű�����:��qR��09�z�#ES:9�}���N+��ΨsV	n��Q�X�E�2AN�![�B���Qc���X[@��'y��\F�~�xK�sb�Y1#��A�=����W��*n�(�R�n�)b�*�e���K���$���0�+u�.!��-@�`E�1��=��mA|(u	��鸢��.]]c5���C� �P��B�5>};[aGvZ��O7F����Ȥ�O��w�eCӳ��(��L�PМt���egh���9A~���������dX��Kҋ��Q%A�b?Y̙M�N�93���������j�G�U ����H�X+�=/C,bp��SsZ����>���7O��	K�^6Gf�k�nͽ�wYl���̼�
��[
 ����,u�;V��s�j@=�R[/2hb�md���kU�Z����g�����Ϊ�Yg��a�W�dNU�*������o�|�uC
�u $5>e�y\��#7��9�]D�C�&��	5'.kO��2��ga�	s�%�i4��=�Rc�tRj�1�.5|q��V!Į�*���
	���e�}׬M�6Rr��5C��ϻ ����Q�kE�
ϼŪ�����mE7ӮYz�M��S<�c��G��)j�)�B���*��S+�֪�{?<��U��K�0ʄ{v����Խ�;
�T���7��ừt���jfs�&;�Y[���?q2Q���1e��]K��-3P�f��c`��!�i,u7�������{3��b��Ƨ����y��Gr\��55��uVqЫ�|L��.�h���rW3���w+�84PP�j�'�'�he������o��e�8�\]��I�.�DԪ�Yj���3g�֤�H���Cn���.t"�B��
Q�
��g�`��M��:�dvb������Ľ��_0������������ I��^����	�&��_���W��1��az�5G�0�Rt���Zw��J�	��9U�:�438������j˂�����K�޴�q�V�u�A	y:�H����Îl�zdU�B��������Z]���OU@Yo^B"�b�l;e@�U �e����� ���8��:�m9T:`9������x5wٲ�͈j����<����ೝ��W�R7c�ݳ��{�!=���#��z�o���aB��84�E|,G�^��3��h�I��"���w:S�g���s�@�ϐ�)�4�aC��g��&+,☱�MzW=��w[�g���z0�x���c]�n2�t�Dfn6z���9�|�.��Ky�||�6��
ӑ{�P/bSYr�+�8P�l��0�lW�Ԗ��҂NCͷp�+@�w�20�+)�A��%�XX��f0۵�4��m�}�F������� ��X� _y�B	_҈�ڙ��?I1�������P<ԥ�� ��3�|k��am7;RR���K�H�B˒U��#�������l�
X8q����U��UsflSP�����?S�@�W��_�^9@�ξ�X�a����,)�B��XLgs\�:꿦3$%Ld�C�r���,w��&d@��w*k���������$�wE��Ԋ�+`���6 &o� �N˄}<���6��k="Y`� 29�r�Kﬔ���Z�|\���-Nx�r�֢��rvV�[�+{8iQX1l`]��<��� �u^������؟�	9 6?�u�+�
�'�O��$P��D�Y�X��'gN�M}�(�H�'�(E���K��ٚ1u��d"�a�/����'�E��#�%E� 8eL'ʪD����ϫ� ��@v1B5�K����~E]Ed�G�hew)S��i�{K�F�XF~�L�Iqپ���4.FIwVm���w��h~�F;��2�KUȁ,6L�3�Ō҇W3J7�O9���$�"k� d���'`>5��S�dӾS%ZȐ���05&��u�j,�b�`;YL�|��!�)��v�b95Dϭ�؅ǅ�L7 ���=1E����^�gCŸ���U0;g��a���dA�E}�K�c���]�*�XJ�1��߷���Ţ���r�s�W/��J�?��b�M6��C�gj-:�@�p�-WU/�U�ѝݮ>�I���w��(Sl8O7������ї�k�o6�CK��Υ��"�$؝1q�Qk��v*6ȴd��?ě4W���/�����$f�í-�,��*Z���9t�nW%$�<�F�o�y1S�) Oٓ@�7 1QR*@�p�q�;�uu{,ԧNX[$�\�n�N%�P:*�(`��+�"�Xn�<�Y�V~��Is��kM����fd��6� W�H�\�.j�l���k��B�>����mב�B��Ǟ�*xuL�q�8��UF�Ua��W�r]Q����_·l{iE�]����-�8"�J(�o�H~g��	�ح0��s(�6�o8���QD���+��&�Y� )sJ��p�5���%"�t���]��㫣�������}��RO|R�Ӗ�ŋ�ck��y�s�Ss<ݷrϝ����v�Iٻň��G�ZH!'�ڙ����j�ց�T���N~�*���s�I�5��̘m��$7E����O��4mÇ��D�~<"�^��@r�`(�i��Z�C�q��
Q�T�~�\�t_�R�Sz��~�yhEfIЂ �'��e���*K�l~�f����y��q;�]��b�b?]�;�7q ZD)R{����vXȑ�����+~����7d�h�q��1p�9�d��g��/O,E��EV�]������o#&���	ﯥD���s5Inlė[�Ņ�:���*#�a/�����+QwP8� !�?ѽ�$x�5�5&>>�h�~�Fk�'�7����(����x-v9*-�Ȍ5ʽ�^��l@�I�'�j_ r��et����E)\��=��,��<�C^�����j�~ZyѸ$/��F<�����LS���v�{��y�q�� +KA�I6~=<�t	Qd	9�a7��!+��]cx,��f�a�DS�J��M�v�ڴ5�_%�ǀ�1܏I�ޗ�l�>����B`?c	���?h�k)�>�}�P��T�Yo@-d���vd=�Ͼ��K�s�#���~2�s4��EC�e�]w���L`���u<2���j�7�Ep�A��{Z����>8�����Q��&��S���}�'k���֩ǥ%��i�d�8z@��BϳH���
�k���^x���6ԓ{��U,,|Io�o�幨6DG-��Y�aX�|t��ѭ��cY��B�Vl-ѓk�}|��v�&[�<�s�Zʵ���Ԭ����9f�uU4I��N�F��g��
1��:��&* Y�&�7K�z�߳����d���@}���D��d��Phэ�J���jz��?`(;�4�1��%���ݻ�y5�����A������ޚ��K�'W�.��.�������J�����$U�r|=4��"����T����M�Y8����@ZE���f�P�В��(�,}��Vr��p�n�5��\D"� �����Z�J;�d�{`����O�e��8�-�͆���=��	m%+O'����<����!>���4��kk\���pG{d��5b�d�Mg���2�}��C�̠�k)��a���%���H�а΄{o߻���n��xa�?�/!�jJ�#8�:��� E�q��!��Q��å�B0�A/Y�a-��j@k�(��W�����֣k� '��,���!�vyC&��TwI�)v��Y���ol|���[��&�w���?e=�V��j�!z4< Q��P�`&��~dݓ/�1�_ �цh�W�����h�D��O�H�����;�}����p�zn��	V���G��Q����?3��F��o������dr{��ɓd�c���{/ٯy��0Ĺ���/����]*������!M������׻/��#3ҷs���O�Y�8[�*��v��^��� W�ܴZ-�e��������]��Ǘ��4��6S����9H#��Z}x#��r�zy�=*L2���C׌aA�<���Gf����~F�	 rX��������U����t^,j�z��x�B"�?��L .=#J/"4�1������c�>!H���=<C�D/\Έ�翰6(g��#D��ԋ'LAC?�s���3E��HX�O���5|y�c3��~�WIJ���3��mvμ;2��U� �^e��_׽�aK�6	9|��FƯ��c�Tk�R�QiM��#)���#��{�[��;x�%@:u�0����+L�N�����D`���(fl{���MA$j����kN΁:3ސP|��L�v�uW�Ԃ��$���jH�f�Y
�!��Y�,)J���b�q��Da�;�%#|�N�Q��?�Y1�g@��4m��P_6L�"w���JTi�(���ɱ]U��M3|ѓ7D���2�c�i��"Nʰa�V��$�oyw�?�M��0���v��q}� e�g�i��"�K��6�x��]�����L�0��~�m���0'��ˏ�����~|Ią -����--���,xV��P�*��ʙc�o��z��N��I�5~H�҇�7�C�3�3�x�������d@407,�#)�}����!��$n��[}B��6݁��J�����HRF�D�g��$2��s��O�d���=zZT�s+5�A�-a�);9���M��[t�1��D`y����g\TI�_�90��&V�K�oUb�v�ݠ�0��!�W+��ys	�8O��:8��E1c9)n����&c#?ub�N>=m���ɺ��?��%��wl�۾�?=��L/��'W-�������Y�h�i�ݤ&���>�8�A�)d��Fb�Z���J�������Ԁ�w�n���I�~
��-�+��(��n��Ԙ�c��2�:[��i�j��z�����o�p�d]X����Kz��|T�d�[1*�Þk5Hq*�*F�MF�%U%��j;����`8�9ui^�~ ?�߱�"_+7Q�y�2�b !���^|ˁH�i�➂Pg��8@���4��J�i��;��M�t��D���"vYw��Kz�Fץ�	{�>��Bwc��,{�ׄux9f�w�D���y���v��nS�����	oU�<a&�91�%�4�Q���q��A ��F�k�}��Na�J�i�3w�p}d�J�����V� }2�A�P�R��ҷ���84}wI�"8 
.���J�^���	�(&hR�-ST\/~��.�d܎���H�b��&�]�M�)�i����L��f��h';EU��*>x�������a�}�)��X�+�fj	���	���!�����P�a^�W�}k���9mF��� &uP+�gt���,���|��s !H&�m�r�zr���~lHѨ�>r���>�d{\0��ph֟q���0S����~�^P��D����֡P�T��Q�80y3���Bgo���12O��@7%���!�oޅ�`�u�Л	)�<���wg���;Kε��sVJ��|�Ԡ�4�Z����dϭ���(x�QBu�6w�@{��D�=ZK�`���\v�ԡ-7V��9�p�{�5���~F�<.����\����~�|�o���Q}!�X[ �aS��K%�%������+�Ͻ�B���I���83�*�
;����%�4���y�b�� �PuQB��1���I�����V@�0�}�� ����5�rWT�i���r1��̎I��A�
8��>���a,�; �`����˪���_�j�w� ��<�F�Q����q���4����Oy^DL�\���+j%��n�3`!R��'r���Z����@�QU���K��}�s߀�M�&T��' �����E�[�f���jL���	H�����b�(�ǋ1[�`0v:��Y�%�/<X����l����������[�ƶ��]*H�,�ݥ���2��B6,�ӠF�qC��l5�E��ÿ�~E�B�$�Ҟr��Vg�'s!�s\���O��5�T�<�0�:ߦ��ُ;�����9��C�e����JV��.���?�Ӓ\E[�d��+/��d����u��L�7S%h�b���՜E�����2Ms�e�����I��$�H��Ok�@�Qϐ�̠�܍J�V���6�+��Y4��P��@4B褒}Cҋ��,���Q��,����b/�ߊ���q���B����$��J/s����=:8��E;��g�	����D���.��b�(�*J��p{�� ����z����p�Qq�'���Q���{��K�xۥ�<����������� [	�4�Ȕ$NJd�6�Y�]u��Y�Q�;��5���駗f)�f����ң��d��0�
$"K��=ߗ7=oFrݞ(/m�o�F�S���X;06��/��Iz��~��6jH��t��;A�&f���g��D��l��N��A�i/hqF�P6���3������]|�����|$3�}&���m�ٴc�M�r���9�:���D���p�}I��W�� ���>�o�ͽ[J%w��F@�������ׄ�k��v���Q2��"�n5E�D����ru���O?7�BKv�0�bo`Ћ+�V%Gm�;��32����P�N�]m�I{\�e_eٸ���⋈����O��wm3&M�	�[�t �o)��`U���'ʸ���_p�0�,�������Խ���d./��/r�@5QF���op�;�d��$A����w~�昿����ȚM�AkO��l��H�4
����2���^-�0NJSs��H��Hz�he���r��b�N�H�mP)�b�2��BU�5M���`!��箝���S��""�2�#y9�Ҥ�1ۜX�כ�u�������[�)�������d�[M�Ļ�'I����`�PZ�]�3�.��1�H82F����H�#�Xj�f-U'�ǼD-�?&l\��>�/"��laS�d]O1�Aa�c�H��B���]�?��qjڮ�
̕����)�4�kʴ�`˔_�2�!�귷cj�j,�	�`�d��QHI5�g���(��Q	����H�m�+.8j�a6�eX�A[��W�.�u&y3��
N�.ʞ`l�8�"V�j�H�+
/(9� �d����?\]�G��?�����<�/�H�Q�f)/�a�c�0h-�ܟ=�.{�n[gH��
V���ش5І�!��h7��_����$z���~��Mڨ��7xio�W��,�t���m�2�J�V�W� �tԁ.(_ew���?�5Qh
X�����{�5��ň:i_ �B�r����!��M���2tm􀵶�n CN��v��.�F�NZ���|7��{�戟��RY:���	T��R�C��M�O�>~��Ӈ��G��v<����Rk�$�Z�ci�?�!�<����Dw�C�-$yL����1�V�Q�7�{�^�}a��ﾭjpm7�SW��� ��ŭ�0݄�4ғdU���7}"�lj�lb����Fm�FP,��YZ�fck�_ɼ�H�;��, ���ǩ�=�m�-�@
�ֺ~u
�`oe�$�w��_��t�.��|�7,jN�f��6]�=ɇ{�,B�Bءv�1G����$L����6��=S�e.������^�휚�Y��Kda�%B�0b��5��x9�`V��4�p�=s�K�BT(�����V�|$W���?���+�5Kݲ��>Ƃ��ξX�F��|S�kU��g�6�>��:G}_���v̔|W�b���g��)��w��2=yȔ�!��}�(�?D��}�s����c��6��Z�\>�����w����m���8�ܳ.MV@��euN��,�{Q��(!?�*.��L,���Ɗ�����\#.���Tƙ�Ӵ>��&��؈! �(7�q?��8�w+�G��wS��\�;m������e���?P�n��m����a
���l{?�c�{�
��7J�����o�w��l=ŧ�ۨ�2de`bʉ��~H�fש�z�d��t�ގr�2���g)��t`v��sVA�D�����͛�X;{��FR���҂�Z	Ԃx�b ��(U�H���e�b,TR'��{���J]֣�<|�g� 'ޭ��Ʀr��~�^�kp��1F¥)��|��6����o���2ף�!� ��n�S� ��B`������}��ե'��נ�MؓO��t/*`(����>�s�q������*�]Voh�~�P��PgV�J���Hmk%��GB�m�N�Sj_Ju�7�|��Ĳ�Te�+���R+8�}�q�fv
#�!yV��ދ���x�J���F=~�@�	�s��a �|}��m�ϥ�R�0dD���1�d���h澌Z46#U�u��W��Q�qV�ۖ���}�τ�r��>�U�0x�޲�R�^�Ǖ�Ac��qc9�����	ğ�@Y���JNEU���/yx�j���Rl���v+���!��� nT�ce���}�!ݚ.���@��\�"��l�ǆQVx ��KS��n|����Q��wh׃�����E�|��}w[92�+B%��A^�ϘrE"I��'k�+Sɞ��>������Q�M~ϥy�;���t�"��������M����7����ᚅ<�_�j
�ǯaq��\J�|��_u���."����>���cɟ��gv8>�5�J������M��ۚ��`4+�e�����$��>�t��Q%�Α���ު��_��Q+�:3 �s8��<�ZGڍ�''�2V��󽶻K9i������%��!�P����:>=m��>�u��3��S�|h�&��̽z�ǉ(�C���#zv��%�֧"L�W$<|Vp�^����ֲ�_>�V���W+O/�.�~'�6s�&�_$K����X�Lꀓ�lvRB!�<.m�A��=����'IKp��*����U �9��#�\p����@~]��k\oOKs搢�t��T����pN��'F�Gg*�{�uh`8�e:���)��������|F=T���]R<3��I����:��c5p�󶬨h��~���U�iH���Zm�S.�Ȭ�)��c��U:�*�:1֚�۞���x-̡j���/<C��Ѹ2���5��S{Ӏ��4��Aa@j�A	����$F��jBH7ΐ�7I�J�f��N|���=|+�?�����A�I��HM3�����B����˥n�c
u6��t�v�ϲB�u�%4��W̈�%��=iڤ�Sj�+�?V^�� �^0��r�����s�Y��cX>���w�˩�H*^S��u޼�ЈϿ:� 4�M������^V��)������K�*�	F�]�k�u�S�G�v��3]��YYr~rM�g?�<TU`�-�U�W�
��1�1"��T��~�9Q�-9|�9�^����x^"���=��FVR�떊��߿+x(�,m�.�[<��[?!��$��u�i�Xj3���H(`3�C�T����a��/��o����hD(�mZ����_�# ��6��Ď/������X��1;�cY+�'�̱j����b����k:{����K8ҏI�Q<��r�b�A3��T�10Q�d�����∊��N�H{������w�P)#��:t̏V�]æ���0�?���7��޻�t�oA� �i�MF���iœ��]�e��q�y
��{K1�,0[�'?,T���~�ST����XcB�"��Щ��rېV���a �V:�@|�Z�W1�k^T'Y3�" ��Ҝ4ł�A�
�p��69��R0��0�����D���yC���	����5��<�6:��<�&L��C)��V^e�nY��Yq�j�E�?	�<QY��Z&拪���FɝQ/���T����*����H5>͜��w���Ga�@F����=̧�)��5�W�kl���o�摍{P�'���]h<�	�%��J�	�C��^.�E!�o�tz��sOZ�f�bHO��P���Fm��4l��&�(q��_�͒<�4du9ӡ:1�0���ic�Q����S1�<?��m����j1V�}�����.S������z;�5Y�2��4�E��ex�d�⾨� ��d2�
��~�q?�q�l�f>T}a�$.�t�]�y�����{�b�A��rż� ;~�9�#ڷ�S��Ԟx.�^�ŭb��]��ej�t���q,&�%�����^ 5uP�l��3n.��x�L�o����(x��1�܀����`�BR��-�4{kbY�܌�Y�I�����^��)&�V� �Y�֡�tΚܱ�[���sfdI;��5��~>n��������
�I%@��n��)�(���H��Z�C"�'woxG�8�՞��VuV
�7��6\G�63�kjcK7ַ֦I��)�?}$�<�d�{J/����&ܝ:�;E�p�)_����e��2�*�X�.l5!�<]N���%p�S4�[�Ȭ�?M�Hҵ�ٲϹpa��l����`k����;�E�q7Q};V�	�%%L���Jʴ>��-t��뵉m�����|��(�����T\bE��b_i�M<(  3ʖY<�Sv�ײH���*�=Wf��FU��@�d�l��j�ld����!D�Ğ}������dr*�ؙ�lBr���p��6EO����b�Tn-�6iɶi+*2+r�2:����}�����0g�?��DGֈڭۍ�`��1�a��Cj��?�zv>|�^��� ��\��Ig��1)�{9�j�/�I�Pi�fd�'W��5�p��Z�������i_֟8���=�A!�d��
�YY���u�	t���!��hK�����6y-�>��OBk��B��%�K�x%􃎵BߨX�	QnU�����:�#��
%�<�[���9��y1�_�����P�>!�ڳC-_�kp����gl?�s��a�.���c"A�weCi|�N��I34"�\ʢ�{�=~�G�r����^bx�����e+�I ޙ9p`�v��T�lf蠎�r̩v!�F	���� �c]uu�;���j���#���j�Q��jZ/mUZ���������7J�U2���M;����Ǎn��nI�@��*~L�^�;��խa���u	4)�`�!a%"�!
�L��Ӌ+?����7�O2cxjIxӾ@��_�jr�����Y��
�B��i�٭��K����7�#~�β�NiW?Y��J.ŻBP���EcՈI�.��\_�&�ZߍeԎ��>ϫ�����+q�E� �(t�␥3������p[&��q�ߋ|���6�n/Ç�ݮ!��∼��(&�f0�}G�҉�\u�!hW�ƄCk���9'��j`1�o��Q�ϒ�M�@|�p�3���\C����=�n�pאJD�3T�)3��2k-hs�~�K�o��EF/D-�^0�j'��O+jͧ;�����޵��"ҹ�P�)c&$��+)LR
K ��(��|��&��(�^#o��h�R#�']K��OI)#�D+3-/�����PVJZ��O)�NBxC2��{�����7bm.2N�{�i�1���U& ���p�9��Bc<�+k/e&��0Z�
�K���0�ij"`&�Rf����t}d���Kicl��W�,j��Pf�{�*�)���X�Z2�ڒ��4����iZğ��Q�[�������;���A���J6���$6�����_��J2T�!��<�u8h>@���;�Y���(pF��0���N�*�L��vǌ�Ͽs֟|�Y�a�Y]�U
�<,`׎y��@
��O�����F���[`�m��=_�/o.�#������OX��D�ͳ�wz�<��	�{վY�O~[\LR��Zo��2�бC����UODk�a��^�%,�{S�:�h�d�&���R�<���`�-9.�]I���U��`��)d���ڐu?P �پ5X\�Q@����w�Oe��
�T?�k�;RC�W���Z��cSVca����&"�5���U98Bp���ɞ+p�*�g�>�"׭߉Wթ-y~?�	9Rb%���[a-���i���Ĵ"�H�"8��1l"u����º���6nR�;��S�B��L�@��Y0ӹ��$Ȉnv����6tX��C:}��"�#�˶��l<���ՐXI�k��S�,.��+�2n��U�o,���Ct���S�ˇ�b� �x���e�Z{�pU_x�q���<��h�� �m�����T��f�f>��tg�~՛E�]���c���ԟ��;�_n�=��p8����2���GM�A�(Xe����|�Y���#9��K%��J>9�{��Y�i�ހ�m��5+��Y��܇-�%�E
�Y�iK&Q[��%(X�X^Mˋ�x��H	�J�K�P�]����b$Av,�j`$^��qNX(^�E�{%m��D��r�����V����k�K=�S＞ku���~�a_O��w7T'ԱI�?�![���Y�`ZW7me��ֿl�G.Id��x���	�-B*�| ĝ�l��`���|���	��e�?x+����Ⅿ*�t�d0طd{M�z�N!u��Itss���}Ա<*�ٳ��j�w��4*�\6�Qӊ!�Q��R�,d7��0q-+U��T3���+�[�
�J�|.TL���b�B�LW���~ҭ؀ ��ȡY��w���3��.U�pTg&�ؖq0�̡Gx��،�Z�#�L�?�^QO�����T�\�K��%�̅��ZO��Bp�&k.a�!��x��� �P�IM�N�*�3u��y�l4Z�r�F�
�n�-����ѡ��1r_�����HN�R�	��Nr�?�T�d.�m-,���� ]�.����}��|:fϩ'ģ���7 ��w�3�"�YN��<u�}9�ؙd(�=�;�Sv��S����U�L��o����RH�K�bb`���^�jO4s�v�yJp�@��Ѧm�%d�\���Q^ố\������B���GbX�
)��֠h���'N�A��琵�8B�1���S����fo��)f���r+��a�5��f�RP�D���t���(tʔ�n�sCn�?Es���	���������d�%s���`��!�`�6Xr�I���d�Pt��4�;�H�i1^Ỗ#&v�w���$�Q�۞�h�*_LgG!t��Ʊ��'��4���-�xJ/6�0��>�D��}��W>�ъ��J΅A<N�@����p�wOt��v��g+`(����\�P��Á��2���u�
�5�ڐ3���O�[�9}T^Z�z�p�vm�,s�Z_[��yΝ�n~!�qJ_)(q)�m�����p�
u݈���ɏ�,��"�������/w#_����b�YW:�Þd�/��F�9Ψ�r����p[N�LD�qU�u��{o�5��ܑ�R�:��U>791G���=a���	TLj�q	�S�hD�_yǬCi��д��Y/�Œ�)���r:���?����3��6oZT
���o5��J��O�t3վ�։��,�lL��1���Ҕ�"!_�D?d��/`���g��83��-���LbY���Ñ����"0�(�'�d�8�kC�1�̌��e�$�?��"O��Ƙa�����`�Uk����W	��A���׊S��������LO��w_y���	�<����������͞{��h7��\dݔ���:�-o����AL���kJr��>`"���{d���G����,��{�����)$)�P�5!�*'kxtr��4���x5�|��E۬��o�Ϲm�nf���#c����ej�o]�9{�=m�C���d��i�;٠I���;��G$N�v�����4�%WD�]ftI��攏F	-���k�9q�.���A��8�(����#��\���[�ԐKb�>�ϓwL� S�V� nXB�p�6aJ����� �[l�븷�g��s��R�|{��y��3<�V�Z<��LXn�*c����pT��Z��*��<PdZ/�Bx����7SeE�@HdTm'NԄ��-:y���SF�3\�S��!�?�g.��p���a��g �6'C���I�	x��I��g��t$�|����+A�W6�-��a�w��п[c�޸v|,�~�(�L��^׷r}�C�{.����'�ļ��O���m`w����!p����
CC�0m�b�@�BCt������$Y�_��x����/(}Jh�l}��^%N��0�|��ᖩM�����6�ݗћ��4���V/,]�Y����M(����v,;�z�㇍Y�TD�o�z9��d��^��ӵ�_K������A��u!Mթy|���K�$hA�H��v]�#�! =ZO*W����
I����lZ���wr;Q�X������e���w��Jր��TA\��)fp돂h֝�����N�'Ďw�>7l��p̨_<X깒�I��N<$�V�ct'r�1-cr֢?��5Y���뺊4��֜c�]��Rqt��h���
����6¼<�a'� 'mGZ�9�C�^*�w���# X�YȂ�!	���� ��\��C�5ak��H�P�- )2k��wߍn�u浯�`�n�*��i�ԏћ���.
�/m`&AItaXH�.�蘶-���s��]_�b����4��x�ڸ�P���P�UM[;r�K�qs��u��{����Z�x��f�������Hp��\B���Ӕe�n�>�%X�k��e�\�􆉎%�SU�_�|Y5��S����ٟ,��qBh+6�؂*�{�AÈ�jX4˿��
�:;^"���\����	^�j/~�\S�[&��z��b��ퟷ��h���?�q
bC<m�8��p@��'�p�Bi�(΁��=��e�扡�%�Ec��
3�����g�D���׃&zJ4�F�YoEz�gn��H��L�j������N�w����QH�I ��0���� ��l�Q�Q��cG�?�En�U�A����d�ܧMm�v�0��9��gTyfx�қ�6$��X/ا|�/�����ol�\O��Qb�y�؏�%�zδ
⩂���mKs.���GKn��
�~YI�Z�����P�Υ2%��ŌZ���e����F�u����^��2�) �����텀K�#i���	r_Jr�	�bwM	��k��ۃp�[!���R�C�C�g�q���)�֋+s��/�>����E3��I޲������%��Ýi{�-r�wrr��l�w�c�D]��:�)�ҴN��%3��ۃq���,�����)��s�L؋%���ʰ6Κ��q\w]�D&Cҥ&�*ì#0x���ב�'WPg���������XF�˥é�*oڋq� E#�Y�
 ǑJk"�Tw�f�����	@R���Ag�&" ��(����O
{:)�]m�c[ �l�4�@o�	�]�����)�*�J�`̫�����M�G%�m�����������V�M(�HXx��jL�\�?$�Q����8B���T}>(�)~�uV��G��u�6���HZ(�s�򩗨��݈���:-���iY�|��3)��Ph�atVn}�`Y������^N5wn㺕���>�߻8�P>�(d������l8�Ld:�,K�u��g}x��P6l��ސ���x_�Բ�5ac�W$�jMr�4�8��»I��٣�V�p4��fE�W��[�f!���@�F.@l�a-�ɒ��ĵ/}� c=�ofdD�A;wL��9�0��UN����e�ۿ��X��o�q������3��~���
�E���0��I�5'�G�iX-�d���w�(�-�2��F@M�P��%�5�f`s:2D�~����D ��3]��?A<��[�/�(��/	h��7����s£À�.�s#�uAf
I2(�ᖊ.��'��p	@�#���#u tb$��@[od
e�f)����J>y&�6s�q��m�j>�;�lhhL�!�p/��o(�b�v ����p����[������if�چ��p�>��載-�c>�-�Xծ1�33�Z���jęd�O�:Zc�e��#�@�::��}?�T$�B����J�Z�����J�
Ӵ�u԰R��:|�l��@�h�8�W3/���:�F����0���s����T8ɺ/�<��4�����S�i�>	/ǛcF,|+{��Ke>��!Џh��N���T�����`MPd(��ц�=e��Pjh�␫;j�R�X@�ԑ�	.���L��sMf�(�ޟ���6I���X�c�eI��Up28�Y%r��!4�n��:/�k���9cX�v�=����Џ�y��x�b�)�i^�]��4�5�e���U��y>�R�tL�W8#+�p�{��3�'����k\+�X ��<=�mg�e"T� D����H繩n��i2�2�z�4?jp�a�݂=�[��A��ް1!���-�	�_�xK�@��Z�6k�vW�s���H3�C�ѥukay(M"�/�0�o��������������*Mt�Tb$)��*�x�׹h|��;��R���V��M������9U.� ��B�-Y5`1��3�e�4��E㦄�L$c�ZC����E�98lLǖ�j�l&6
���>�	O�*��҆�X9�|��[[���)
)��F��������!k�Y�5A
ͤ��~ӵ��g,)�YxU]�k�+o
�tU�0/&6V�c���R�,��l)�H"���`���*�n/�?{Dۜ��J�6<F�4�@�kܖM��p#�)R�;��Ga�	���;C֠S��s�Ҍh�E��qWV)" qz���x-,l	'������ԩ�k�]:�,��T�4���4-ᑹm���·_�y�Tjعx3�L�L��y���3Y�K����4�|+�u*�0���+����!*�/��*G��.�2�2�KFc+�V�0MG�H���
`��qg- �625n�tv�_S��ӳ�\����N�J���Gn)���U�e�@�֥��"bq���:�X��&|�i% �ؑ+K������+��	2��@!��*.΋��� S����p�?��L���D$^￉�-�Ydun�~�׈:�k3Q̱rD�O������":sk�`ݶ�����.��w�{x���	<�N��o=/{2����#@2��O�D�p�݋ᴑ���^dLl��G�f�A����7"ȗ+�B��������)���׉���Z�g��A����dOi��$��)��Q��%6%�y��Tz畄�֖�@|wU�.X�0��0�%�9�I��7��-�:���P�k��]���W_�O�Yn\�RU�^W�܈7\�"}� ���Օ�u� :�M���{���S�ϝ��Z:��	l4=ɖ^q�}�V9�ݕ���@t��֢�R�*���l�1�IQ2�2�P� ����>� K�6�ǒ2RϘ�J�6z����|բ��hg]�i$=��2&X�7O��9?~6v6��n�I�p�"�<��Oۤ	���m ��?T�U�;M�F���E8Ȟ�x�p*�7�g@�5�Q�[��\�Eb���"�9�K���R�+�%����	+�YB�hM>�d��+@?gd,]M�h�B�t���M����5$����!@$��P5���O��0���򼢫�Ȳ�g�+�;+�H��7R�0ǭ���`J�\蹐��Xj�*VMi+@l��,}PQf�A��'����TM��V��K�>~Ms��������~�����4n<���������	� J����Z[�V��<>�D�^�>����Y?�bc&Y�l�D�a��i�P{(�òN���̠��lJ��=�e�E��EI������#T�+��Z)�&�5�ٺ�`Dڞ䚦��n��ɸ+xT��-��=߶�.�VK���]�A*������<5n����k�Q[����_*��w7�R�����N�9;4F]G���
X%��2�[��_^����_����͏��IUw;���h�dY�6C���U�*�]��kiQ����#�r�J�>�!��Ak��f���m�F�.��̄�8�;�4���-(Y6�ı#.��� ������AsR���u~%haq>"� ���%���B-I`Pfk�y�b�a]
,����;Z��=��z@	�M������e�+�:8-t���f�\ȗ7����i
�{�c���[@a/D���l�ƴ!�WzT!f�E�i�ϵ �=b��0n�׶X���FP16����L��ۭ�~,\�����PZ/-H{i�"�{��q�a�8�]��f�4���ŝr�Jm��FÓ��5����)nDA!C)E I�T��z��������G��ri���>�:)M�Od#PV9�J0�@A��} 4{>�bԀg�a�,�/u�m����Z� =�-�|��^���50 ����b��Ɏ㊘hȎKD?��{H�K�����o=����� 6G���=}_������f%\ěS^�;;� @��*E��_m�RB����0�mʅ��ʼDIJ8��}+�%k�2�}#��	�JTC�Ѝ�V�d�q�0Q��5��q�`g���w}����Q�I�p�Ϥ?l�
!�Tb,3��
��b��TE9�Dn�b���zuU����������D��@�6R5�
��)k�f+UH���=aX�g�&f�}|����̟��68'�5W��-ҫC?����lD濂��%h}]q�����r/E�����m>��N��*Дs�_��ֈ6tA	�(e�+p�y�fk���_������'�)�w|�xGk%�,���Fg/���,��4�-�t!��{�#�#�{[��R����.��-�W?�<I�~�a�)�'�Q��R�,�K'ׄAiƁ쩃qDud7zJ�'<��no�oL����/��:��V3)�Bq�x��J�0 ��^,��ϝ/���{1��>+�j�)<���'݉8�����ڦ�>{����>3���]K �T������/����Q�������Y�$ �X�;w�K9�����޺�m}v >�,��.�I�%%�R8�jY>�O��N,Gɟ!"c7S�oEw3:�lD��{��쭆��P-�X��ɲ�U�,��Z(�~�Yj�,�MX��F [ڜؠ3�h "tV�`��w��~'�W��|����W吚[$�������������`ÓE�$VC&��Mv���y�+�G����/!3h)u�=�G���2�N�ı�oS�>��xcy��9�� 2�Ҫ����1&�ml��� "��4<�(���?6��[P���7@�w��rI_l' "���l� ��`qq�"��L�Dm�v/�w�!���SF%��K/_C�?{RP�-�Hŉ�%���!�]S$P�����(��B{`�+���֫�{IsGY����Þ�L�R@��iV��!
�œ �2'@?��=�vK�N�9���r9�̀?hZ�Nk4@��p��N#v���8��|���N���H[U�(F��r��/��̈k�Q����J�� .�'�,b	)j~�� l�}��aF�j�E��)���Ø5yzNi�N�E��Ҏ�(�� wG��c��?��$�s, l��I�nO��/VjA��;alU�\�m/CG�9�)v�+�O<M��9�Yӿ��,�R-$F&8��" k���M�BaN��r��S��u	��5L3���&��/��{l���!ٸ��8���0��h�qC�\�h��se�4�n#VI[��q��ףU�Ϧ
�鏱�
���&�W7%7�!߶	w"ݼt��F��E�~(Q�� oZI�PMc'�%������jc���Ⲃ����^�X����_y�|�M���]W���
F8��~\�k�HH�8���䘆��NzH�AՀ � �엠�X��=�'���ᡣ���������U���}����(�i̤���%�w]��Ñ���-I�9�:�w�sV哥�E׎��_��k�x�g��
�������`Z-u1C�u��Na<^	�l���!㨼L���ed5��B����5X��\����Lr��r�rk���`�#?��wg����Ŷ��=E2t�O���o�%3Π�,ԛ��F�5��>��4糑����,�l���k㻠C�� �Wf�8^G��Ϊ�>��օ�J��:�p��?+lK����2m��g/e�~kCsp���@��Z����hy�ٜwy���4�h�4֤w(b�D�E��Qh/��C;�6D����#�v�5�Le���~���{��?�͇�-�*ur�8��B]��xv����˷Sd���R
�(ZV����z��c�&���H����Ȣ�г4�ll������ǵ~M�}�'�aG*��*��i0��Y�ژ8%�B�rY�����\�<�����-yNf������S����_�}�T�໠�> ��~d�,�GL�ŀV`ȇh�Ұ�+$��ڜ���'�Ma�G��E
�DySO}!���:Җ���l%%� 	䠐:�O�>Sӂ�X���W+'i��{�d��3��6��/�7˶h�kf9`y�Wď��
+TH8g�?䵭���$:�*q�=��ȓfo��?�|kBC��<�&H�ZUH��]��Xg�E_��pO�b���(pI��;�=e��_�����;_��!�G�+�-S���V��{�=P�@0�߶�����d�9Q��GF���J��Cn���x�䜡Y싛z�g_>�u%�	��x=o�;���~���D������zx�X�lĴ$IП��;�W��(dl=^�����K�*��]� @O\����vc�5��n�x�WEY���mC��alg��Z��?�e�ơ{��h)�.�����%��*�.��Ѳ,~4��uD��RE+�v�*©]��q�����o�3r�8B�Μ��	�P``L�m{j��r�ik������*Nl�LK�)��Va�(���DbU�����/S�x%y��9C/hw� �Heh7&�A���	c=��a����3-�i�>�0�����~(�Y=d���wtԉ$J�w�uU*A��#H�{&�v������Ǔ�M�-`�N݆����\�(X3�
�)��ߤ�םМ��ON�c'\wrk4��!Z��E~� ��9�:�U}����<~�\�ryx:�b�.!&�~//2�H�o:O}�Q���c[b����P%�ipޕ^֒��խ�R�|k�P.��KԊS��H�r�Q�}q�R��k�cc]����W��U��L����He��OP |�O~��hc�l���N��5v":�V�S�.�*�� ����F���JwW�]'Gl�呠�d�<���K��QS*��8
wYG˰̷�	U7�F+i�kTPI�����S��\��?�}�e1����:�
�7��m~*dE9z5��H�w,Bj}8@��-����@�H���s7lad��9�g-ح5CɜcTe)7i��n���;����>�黷�>��Ժ�Dl���çQ�b;ܶ@=���}�`�i���iTN�ǟ)y�#�<�������C 5����I�tL�M|��p���[!B��@�u�Ƭy�M��Gg��l@JJ"'��8�c�`v���cgZ��L��{�Ar�۰�k���%�'��o�=��%M�M6�W����p���;��r��%�TCmrb��Fgp-2����ʧr)^�HX��LwN9�ɇ`�"Z$#."�>,�^�w9�� �߂��܋��=��4�]�q��o�}��0�4(���v[��v�M�]ɊK;n�
`F��sD�����x�1p�L&A�O��@��<0i-ǰ]OM�I�@��>J�GSX��w�l�g�Fk7dB�o؇�j� �OV�y�k�����F���&���h�^��o�ֺd`o7�Bd+��/\�)ʵ��B�[Q<�2-.���g|X���r��ԯ��4;�0�
i_�X���{����Y�F�.c2\�]���ѷg.�>��c����\ S�[N�����m��0<Us�]烜�����Q��3qʯ-���ӺաY�4W�G�� d^ʤ:�h �,ϛ�-��g���6�nP�� ��\P���_�;��,��Ruv(ٿ#u���=�}.���W|/�MU�iC����|4�����U^�MC���A��ΰ��:W6B6��`�W��9���8���j
���s�����c��G*��F��y�Ǟ�N��qu�PJ�JA��*j�t��U��gEFY�(<d߃,:�듎����CR���
[]⽪ZO���g�D��r��Z��X��WSdm7�r��.Ij����=N#����=3I�R��J�:������nK��y+����q�e\��<?e�J�^�;����ک*��}��
%&�)/m��v��u�r�rK׺�oݔ��#�����!�/�)|��+qq��	#
W�C���Np�p��ߟL"*�X���5�p��%3!@�����:�j��E�c(��+|���g�}�f��"0��!úr�#���«Ð�G�u
�T�݉��Ȓ8�9��ܾ�V�H7�~��W�2��{�0�P�$���K�{���P�hՀ�v@��X�U���c+sp��;�D�l��F�i���"Fv`y�\���`�Nl�yYo�*����G����xH��A�r�C�mY%�w!�B_�����=_�5�=0�q�G�E��&�� 2ì�g��X�l�iK��d�A�H�����耩�g"o��Jrw!�xE?|j��\'2eȽ��OB���G��̩�4��G���w����ϧ�,~˳�����b�_��2��7���^Q�r���Ո�Ho��Dy��|�2��6x��CJ�����UXPdϦgZ�Gq�*S��ϵ1	��^�YI��xQ�%q�Y���'cύє��-A�,��*�Cw0��⟟�Qb8�Ҵ�TH �P�o��Ћ`65⇝H�M߄U�Q��;i����W����pA���G'����M������d�R������*O���j���X]��joK!k�[]V)�ݓ@��\5n�j	jg�@�[4�(	�ź�b�]d�����6J�?���PqM���@A ��e � ޘ������H6E�YM�b}�i�YmNQg�oi߁Nf��n�o�Bةa�g�'iU>y���ԥȐٳ����G�#�b��𽷕$��:�D� %R��_3��U]�KRk31(a�\1�C�w�2��C]����T(x@<M ��/��o'݈�s���B$���)���z@�ǳ��h�,"�a��)	#����d�Ec�υ%�F4B}hڹLQB
)�sS�<P��M��)W��[ְ��>>������Y� s���~��r�gEg�j���o~�o�
ֺ[�c<6j�M�����.g�h�'�<�`�=�B��*�QX�"���Sc���M獪D �7Ǳ��d�SV����nno�?"
a$�`�Õ����+dR�������0����@m9zSnBĘ�`ȐBn5�۵-�ôk��,���u�oG�'x�j�y�����'(3&���G6c����p+�p�h�aLM�4�֑)�KA�:3��ڢ���!��R���5�'���eN�H�w�ߺm�XTζ;��Y��҂�f��6�\��P6��؍S&�@��3����p��գe&S�������0��/]Z
��^������v�[$��XD7��XE`v�/n'��e�[��`&V�y!(K�s|$[pD���8]s�,�&�5`����7������ϙ�9���O'6�|o|g��.�"��!�����-ZO0z��G'+.LX�W�* ��QHqn��D�;h��Q��2�M( a��I��M��&�K0w�qO��UE-h�;�uKz���_�}u����_�N�m�wl�󽡒�M��,�D>u�MTah���Q~tZ��=Hǈ9٘.���`�wW�Aw��m� Ý/rU��Ե |��:і���b��G�.���yBԔ��W�#�z�Ӝ{��F��HyAba����̄]�t��R�����&��5k�ZvQ�+DW{�#���\'%���H���$�/t�����؊������:L����@�O��Ɖ�\4q/�5�� �p;��P��
�	S��9܉�a�-2X�Nٝ.�+K�3x�E1��C���,��h��j�+�,V��	hfz�E�.Ng�����Zuq�7��f�!���Hg���W����`X���0ӫ�|y �f�`�v�b�b�'ݽ�r���{�"�*Vw[��(�"S�9'�����픯���+;��'O]���&ѵ#����~�d�=5����=(��\j�k��?A~6PW�J��.V�Z:ɤ��{f��OI��Y�I��|۞�.7�y�E���2r&�=��)^�"��i�Ƅ�y����NaoO�������kw⮏��k77����*���9vA_�� ��1�8D8bpq�^d`�_b�b�Q���e�R �Z�z�sf�������0
x��`w�{��G��X*dɐ��])��h+b[�5�[Ġ��o���+xo���s��v���gkL��\��q��U˕�"Z3��r�"eU�����"�C[$��ތJ�V�*��~�6����J2�wd�Z< ���n���ቁ`�P�L��3(l�$'y�j�9L<T�/���-�ٝSeg.�4�x��JЂ��C�΃�s�F�P��=mSF�P�3:$� 4��E�Ü���pH�n-�z�
3}�Y;�w����s3���qqwB�=u��ju�!�����&�
V�B��D	a��f}��#]�f7�?���V�st����L���/�p�2;0�$�}�A�^A���-��Vt��NI!��$m���
��>��3)#K��c�q�����DN�nƈ��2����_oy:��Ϥ�\p7���2R8�� g��[�1���B����aɠ�ӭ>��!`}�:��O�>O`R������*{\���	 OKW͕�&ѧ%�TO?��)���Z�`���Rwyğ�OIop��\a@������*�2��h����sq5Y�ޖ�����;������ڔ�:!>'�|�i�A^�+��g�]���LM�딂]8��
gng��:��e�s��l;�i)�%�/Vu5���GX��qH$L��烓�V���jvW8,�`�뫭�]8ۭ\#k�m3�����wj��OuޑMG����m\`��.�:���)1��%@���]��=��a��:T��㸇����Xc�+S-�����.�-C���%���a��:-�n��ݰ�D�q�Y�Sy�#�t`�����W"!wy�_��s�8%]�ug��f:��|�7p��[���#��ԯ�Co�zX�|�,�'�V�>Ɠ=�-���];�w��	H�>�K�\�X��$60~��(L�T/����Kjm���e�^;�����&Uϱa��D` b�#Ž���-�vJ"�h3�q��c��d]���c��5�྆�ȟ�4`�s�J�]&��u#B���bE��6ٟ�4�51�=�R��*Rc�BTs��ֿ|W����?�ū��R�v��a4��+�\d1�(�:Ds�I��4�x��k2̿����	�8�'"t���~��a��t���W`�k,��Z3K��BGx&|OB�T�<"��)�,�D�����t�L��s�4-.�����sOs����+p�{��L��q"9\�Ot��:�G�[�^0?l��4��H琻%:��zE�D"�D�H5s��e�`cՓ7׬�k�W�����\�rll8�^[v�>�Q�LL���*�]h���6l�çQ�eqXQ����=�$���ބw!Y_�k0���}�SJ��L6_t[�*��Ls]�������b�	��A俜;T �m1��e)���;��֔ �Ճwkq!�������?6 mRx(��������6ۆ�$B�ԁ�>2g�gr+~��s�=����_8Nd�O�,MC��)@�C��!p�\��+�;����<@��1q�-�f����2ƿ%m4{�X�`�X2{�콪�0L� w��j����:T��@�C4x`�@,2��K���������e����w#��43��zn1D�OJ�8�f(@��N�ɡ�8�X���+��^m��s}v|'�Q<����Ǔ���[Q��?�N�|�HG`Ȫv|Z���d�2}]p�ǳ��N�N��|���J��󛣾j�a?�wx@$М�q�u�1Q3A���٭`�g���W[�J��"/{�"��F(��ΨKM{I�a�q�#�ߐQ�l�%
���zi��G/[�S�So�J��m2���k�$B\��O�E�8�G߄5�rLxd;��ۤ T*�%�_��Mkk�U���2�v2���Lɻ���Ij�rX�/c����>k�.�?4N/�������G+J����~<f�I��0�xmQ-�ŀ��`�>��o�!�Y���~X�����4Gcyi���I+x��(�v�j���G��[�mZD��)��1��7y�Rn4�����!Ч�C
���|�~�T�Px��*<�U�gt�w�LE���Q_5U����I
c"p9A7�417{�t-��=v����W���D������5�����1����	�67na��R�Q�Y�������ͺ�d�H�|�ia ���r&�?����.�t�@2�N��p㴡��ĞI�ǣ�[��8W=2(�
Óf���cE�]ϔ��h���gk�p 1�Fm<o�ՙ�%�#�Ö��-	�Qϡ�)��uD]_'a���cZ��8E�5ΉD�R����Ի��7[|�It��"�-3c��c����p��I���b���d�lܖ���2p�{����f0_��ih3�V�R�Q���F|���g����u�;��YU�x��W��]!��S�U���)�'̷�:a�B��A?�QՀ1��͊rO�}s	�60>�8f&����>����!y��|���u��:Ɯ�>��|8��$�9��b��jJ�
�m���'����bX�c������pŽ�FoP˿�
L'�"w�)�����n�Y��5g$d �Ha��rӌgz'�;\^�����������,v���0�����(*#!2*��V?���c��[&{�䠐L*7O*�]��@1�c�t�j�;>*/=�/�j�Jy=��9m�ñe4z�4Nn��D�#~8zZ���H�)t?,%�G.KQ�4�9�h 8�c��i�.#͹e��	��t~I��9�o�3�$@D�3ء��P�fa�!�0���F1'���������f�
���i|�^��O��mZ�����bg��!��Q�Wy:�Bv� k�ǔ߶n2a�6E�6��9QN�yMF:߼�X�����qQ*�%��l�-@W��Hp�{�EM����&H�A�ӏ@�s��#2~5����J��HF���y�K�����`��[ -AT'�E�COӎ��RB`j^t�[��a'WZ6��0~r@�zʴ�u��A5��V�*��**tR&"���d�w��U d8!PcD�
���nS�޺�~/k�������Ū�
�	�:i� �]�j<�17$��Ћ��A�V���ENl���A]�[�9[񢀑�e��'H��QլD- "��!�̵�����eD2{˄�(��aŢ~Q-��}���+;�xkG�jU��b�28I�M�3�� ;ſ�4e"��x��e�c����`}���/���4$��1xܾ�6r�"o�l:�*��B��:������	�|l]�%�������d��;  ��[+��F"�0Qc
�6���IX%�C�psGh:�aU\ᴧ�� 30l����X4`B����H�2e��*y�o�q��	�f�EhZ��0ֻ��؂!>�LS:Hp�>�4�!i�_ag.�gUf^�������YzVg���۾�s��}��Ua���w=?%&z)�Qpmrҥ	&[qJ;R��(c3� t��UE��5�p��O��#)3W&�9渔�������Wz�#��{laV-�h���̛X��Q��%oVː�.�����J0�&O�b�i"��\Z��,yI��e!n���U�9)��d�{6���^)�̰W�>�1JaϾ��PZ�V����f�]����S!$�h,
���Yg���w�ShH�c��1�*��ҝ*L�V,�
/�pP��$�fP�Mz����ıc��q��"���E?�[q��%�U١��&����V��a#?D�l���&�o��W7�< ��J�K�ԙӿ��W3�J׏��\��i���u��S���D7�M�F_c�ky��Ƅ�#|t]�G7YA�
{@�4�(N�c�X��l�{nSgi&c_�6�Gd�;�9���5?���ہ�*u5�;�b�
ba�;��nW=���[ܕ�yxi�*B��� Y�_�����^r䘅Mu_����F�I	7b�˙R�F��f�����M`��eN���@��f�l`��ϟkwL���%�.�S�7�s�ۑ��o37���*BDh�E���n�����fi�׷8Os}�[�^6�v�#x��;�c�k3�z{��ױ=�IK�%kE
�xE�\��'v���N�LXj/�Vh�ו'h��םެ�������`{-��8�]�#,�����?�"0�F�g���T���Q�ݒ3
�{�2yf��rK,�PDy�ndhs��V��WP��玹a�օ� q��8���7��4���̱ǋJ���@�
��?!��xy>����<NG�f6(|ߘa�[��(��^�Y�W5� ��:Z[3))��U�H;��C��ͮ�Uw������͌/�#�	��O�;�XA`�-L&��4�L�%����L���ܐ7�����S��J)��fL.��d����|]� ኹ`��k�� e�YA	g\�>#�� �������m�2p�]	�*�3�z(��0�lBӼpK������Ra�|�9�qԆS�I��7�D��熿�/'��A�[2^5^�۞{:0nC�ٚ�������V�Y�ڤI��!�����f�.E\x���Zw�e���<S롁#	21o_f�녱�������N-�(�����������ذ���}�*�kmɟ`_-��aֹٶ�]���^D��xȋ-����#A��yd=^����KǕ����>��U�,���.@���D�M�E%���ڥ_`�G�$Ӛ��	�� �O �����*��)�+ٸ4�o���ث��~<^����]�����*��8Y��.����Aĕ$��s�R�m�Sjg�o���!y�^&�,�pOu����uK��.j�[�;��VYcϟ��r��['�3`��U��{q2�\���}��������f4=�����}�d���Y��>â�z����-|��9���p
�м�[T}i�\|� �	�� ���Y��]˓�*���v�A��ͻ�N���yǑ��v�͟�������;�������碔F��7o]�Q�s\&w�f���*C�Tg��R�������?
 �lm�$R��eS�i��G�W���U�0e��L��s��X.}�_y�JNQkuH�W��A��Uv�<��?��jBi������o�R���f�cG����ȎSEGK��0��,��\�����+. eu~��:& ����Յe:9w�|��nI:J�fԚ��G\|���ҙPq���WI{ׄ/�����+�k6��w�w&x���D�����3��+X=(�4�y�Az�R���L/م�0��
e�6pן�E����ԫ�$��_B�_<��:pǸO�޴�gt��"Od��Z�.��~Я���ڊ))_<W�NLtO��4XXb��~�֫Bt�S`%�q+ e����M�5d$�h.s�m�Rx�D�=�#��N+�^�~%���v��!��+�ro�%?ä�Z�l�h9�]�g~�H3�p���N��Ds��q����+k�\�i���(���?�	A���e��⫇t�ȋm)�_k�+&O0^3
�t��ԃm������(�l��dq�������M櫋�X`�����W�������`0�3�^�T_|pdٖ��m�Z��M����v��R=dJb�Yױ��j���B�I��h5�n-�YWZf��� �us�n񺹞t�&����é�,VE+ɜۡ�h"�.�t[mi� 5G������5;�֟54�?m`��=xS%0��Z�?��u�}
#��4"�lZ��3�_rW.���6����n��A~6��4�|t0[\P�ȩP�S�f��:�yD��e������v��פb�����:���/]���o�����, �ɨ�������B�#>����1?�!�`!,׼]��w5  !�G� I�X<.̬��
zϻk_5��w��+.n׶7}��G�m_��ܫҢ�k��S��[bW#p��+��G�n���/Vx�=���1�P	{��KU��
�&  ��n�ƥ�Ԍ�����DI[�B!H�8��i�8y��'�n]�^�c�A&E����|7%Q�^0\�������]\��C%�ٛ2˶����̮T[>aǴíU�Iz�g���
����B)"L+;~͞�asx{QM"��8P21F*��MX��{��-����2784�(y�fg�J\?��u	@����X'?MO��W���b�f�Ͼ�qZ��D�x��zRO5k~��߲���͙��ޫ$��9~B��d�If���郻�fB �a1�2����{�p��8<S�n	d��	����@�}����K#*��[L�_"��z�h>QQ!��� ����R�~��R̷�,Z/��Y�F�L�-��8�s6^��u&n>�k�6����)({ -��r�E����;#�W�Y,��/���d+pϏ鴔�>i*��v�`jz/Ê:~7��7SA���ذP�4	H]�ժ��e�q�������n�,2kbp��]��@\���B�XEu�L
�h��Z
�-�ӕ��y���p�©��I�I��_V���L���])oU�������:�.4C�����C\��^�o�ZkqT�2H��'��!� ��"K#��n�.˒�}c>�*����^��EfN�ͻ)W��)�9�%E�!�p#v�� t]2���eG�Zq�w�K��^	x]ʳ���1@�-�
(�A�Qt�
������0�f�~�p���:�uT%2��/6Y���`��b�]Hk�b�<��#x�'|��^��%� �2���$&��Z*Y7����Q�&�AryFU��7~X�1�H�K��|
��S�f�b���z�����,�%���U �T��(�e��D^�I�~�G�����e�r�;��;k����=�����G����3��u��q4޳ޖ��\4($��Y�	��hn�B>���qO��_o��&�i~n�௳d;ϒ$�]�>;��嘍λ'��xum��3�d$���w�&y��c�M281�.�E��Gc�?4^�3Xq��/���7��$�|[�Gܡ=�0Q[�%֠�#u`�G�z&�J���l(V!����2��v?c@�������H4�������D"����Zˮ�|mj��U��56`�|��N5uTv2ۛ&	7�����K���|�d�jBH�	����X�x�QA��)�("NW�X�$�>
<f��a�d�ǚAQ�v���W>��sq*(bh��2s����X�����x�7%G������.����#�`:&�k���K��o����~1>tQ��J�ą���ڥMv͝V?W�Cj�,*|���.�^K6�,��2�<�{��	-D��N�$iS�2{�A���G؍C���S�&����R9�iX�N0���7�Z�vp���d�RD������y�;���rʗ��`��;i����a�� ���)uv���ބed-�e��ȋ��k��q�;���N�.Oؓ37ե晱�ĳB$qi�{�_� ʔ��2]�㴞��+�߂��-Īct!^�C���h�����k/�)����ɑ\�G6��Zvғ(sw��'�i�{�=�b���Ŗ�.E�əňpx�<&��S���v����_��;�JN��)��n�SG̶�0�1UC�ԧe.���+�M���S�{��!�^>>��w)="+�ѺB�|Ph<���hp9��Yy���|
��£�۟� lL�(y�ƣ̷���cƺ?�s�D�!:�o�#��#��U 3�6Si��D,�M�r	>��HwU���<_��fQ�Q�C�-?4�9��J��(6j�ס1��_d�'�ϸ_��`�?�$���n��jpH̶����R<�� �=�����	=LT�ʗ�M.(���߯����<�O[mTPgTj� �?���C����#vO�H��I+6 �ku���5�+i� ���m�f!��#:m���w�:��5���z�nC�&���MRBg8������7BV�	vo�W~�;���x�O�ȳ��X°�T��_���{��i(�Y�!��)v:�o)�g�!ϚY��Ū�
����Z�z�38�nV�OP�SZ`L*Q� ~�<����CF^�,�_�v��?�Mo�i d�-S��HW���o1�꣖�!;4*�^���D�C�i�}��YN�\�`�\��>�[�Jk�!iS�E�8�s��X������Ǹ,G��M��Ƨ���{�Io3���ף�����#ēv�A�_�P#E
N�A�"��E�4���}�+���X���������m����<�qJ�՜�-��f�>W�!JPN=V�i*����S�K��
�&y�<kY���s��_\g��9R��SEG\�[�᭨��%�X�[i�AR���'Z�ƀ��i)M}�rb\�W�S~�ލ���ztz���Ҟ&'���4�W�`GZ�t\(n�~1u�}�$3^p&@��t|ׂ׆=XjTُ��@[�-Q����J�PxW��bj+,CP����ҩ ���(g^��7��Ⱥ������M
6�~���v��[=A_�<���8�doZ������P?Ҫ�K���~붛#��L%Y�����M13�3�����Z|��@`��]{n���L�K����������{�Y
�a1��)z�0�b�b&��������V[	ҙ�Z�A	�[]�x��I�|����$ӈ�ܸ�#�Ќ��R��v#<\d�?�1 ܊�|�c�z�K���^D]yԨ#�"���,��뺘V��hԗ��q�>A���]����Ɂ����E<v��;Ϗ� �4�J_7X�^�Y���zu*yw����h���E� ����7�h����j���"�>YO����@cT~j��SS���U�l�
P��w�^&馱���� ?�H"$���p�e��~F�&[�h���\�aڐ�kv�
 �:����a��퀾MYeB^�LK_��a��k?�H�����!A�5�,v��&*(��II�A�u~'��"Ͷ�+�g��J�e��	Ꝉ�(K+BںOyMh2{�)��GfpNX���A�#
?��_���+oy�"N�5�)���>�P8�v�W`*�r�L՝pgAh56!�mmJQ�f�{��|X<����?��3�Q��7 �#�a	���߻X".үNʖ��ϲOHybMc��М������/d��O5v�DD���M̴�ތ���˧���:������ÜQ̾L[b����L4zg����!�[I���~��&�p)�R� �ۘ*�b�,�?�/Ժ�2�v�.�!�2<�ha�Q�n�j�Rq�i�2_>�9���ͱz�P��uu-,wxF��[̮ӿ�̱�w�WC2�wV�P[K���#�Y=��J�O���iz	��~�y��Е�<sCsu�?�+І46kff_]3�d6�ޤ+5����v���u^p9��}��
ѢV�x�p�e�kKس�T�յ��{�3�����&�ހν��F~M�!��,;��\YE5n*������%���B��l��������R"<'^�U�#]-�=c���|���e%em��v*X��q�,*��E�p���"2X�T�P,�*��c��ǟ��z'����a#�W�U5.��.ѕ�O8�j����R���U���������;��4#��������ڌD����l�,u& B|P-4�|p�*����E�����cʓ ��--�r[�"�l�]��@��3��c���7�P�t�d� ��PGV�A���t�M�E�2*[�^>>dX�߲~���W�Z�2��)X ��0�sf
�N�A���S�D��{��	x�kɾP��k��W��bs�\�����I��~�^���d�����#��)<��pҽ�6�\A��m���\��P�h�Ul�WZ�͌ev�>p|�L�b	��D�Ƴo_=�_`wc׭���6wq������Q{~U��r;�6��� �E�OM=��o_��U��r3�����'2��@�]�1(���>�0�������A6@�J�B!z]a���{Dh��̤5��Sފ��Z�HR�ȁ'���.���,r'�~h�t�sI^e�J��֦Uǿ�|<`ޑ��Ca��r�N��\G����I��d�.y�3XVD��>1 X&_�m,T�^-B~X�8��W��|�|�^�"�����6o�M�X.ҿ_�v���7j�|pb����}�=*�PhO�;��i�5t�B�;���q�KK�tF��Hg���1nS��4���`+SY��f4�B���P���p �&���c�7a�ӊ��0el�׮���� ����i�IS��SѴ���Rv��CC�YG7��e.H�Zz��0�^��!��6h/�[�h����[_^��]�C�y� ��������t�Pr��%� 4w�M5�ݑ��P�/d.��.vs(�q��$FrT5j��
�6+)�2�1 D�L�^�q�-�9	�3�ˈh�DIG#ݸ �e�'��!N�Y�W����jNit���,|4GA}��!{c�����T5*(EUْ��nG���cT���D�a��5$���1����BO��#Kb⌉���=��1R��/ F����L��g�yeF�/����Xs���W�c@`�����eM��1���2
Q��:�w�/�}�J��7?<vh�^#b�<k"�ȶ���U�$4I����}y6�j��h��|�E[�Җ��'�e�Z�G�����M����ls�G9\!��9�Y���U��۱a��C���� ]�� w�r����Ir��[s_���h����U�q�%��g+���2��mB�!y4N"�mܛRI��Ƨ(K�6����� EF�*:�
9
̀��F�Aq__����.n�ʲCW1|ه������#������)@W���Q��D��!�^)�:����$�ZD=uz�?V̤��4�[�K���9L��+�����N�k��h�"�����r��Mz	��Ebv}fb��!�L�(�
��V� aR�nMM��֛���e�5��p���W�.��C�[e��o��d��e[տwkM�!�h����,?�� i�dgX���e�ܶ��@/���ֱ6����K�̎�g�Uk֭�-��� >"h���S2Do'f����R���0j���`���.ޑ����x�&�ˏ��,�>an��聼H��+��Fy_�7��y�&A4�쵦�6�������� �$�2�����N�Ik!��K���G�������11��e��<O�P s�4� x�e��40 � �Q�u&�����x���u;Q�|R���sf:�Y�O�f��$~Mn7�-�#�]�}���y�qC��[�AJ�M��{��|T���_gS
-n���\MӾ�?5�2�˦��Ąp6ۿ����K�W���|������#ze�a���<���3}�b8��rHY��^W�������w��>����Զ��+��]�&!�C�̺	aY#����%=UZ���}���i)Ȅ���"5sޟ�dTZ�2v�ȧ�FwH�"9A��*��9�F<aiC.�ARV}�XX�\P��@��~[ؿ�����C��U8�,V�g_�n��/<T�Mϱ�5?�q�OhX�������� H#!��0U��ԫ�K>���.���Şhï'��\A� ���Uv�l��1ظKBh9�����#���WC���n�׾[:r�Zvw�⺼���?L��7������[�p��B`��C��ɔ�p�:NP+�����(;��4�����k9f����Ur���]{�f�w�k��	���)�x�N1���ߊ��FXtHO������V��u[��-�7���G�$c�p�)����DB��	�����Ƙ�{Y�9��ٗ��Ŷз4*9f�2MI3$�L�KÆq���{��X�s��rR���wu�s���4���?Tn"�E��V�y�c7:����E��X	LJ�]=�[�Z˅�P>bTb���fH�!|��Л�y�P��JU��|����0�T#�L��K�`Sl��E�rͧ��B��+_���*yKI�lX.����u9~o��gVM?�f��q��7�1��}�4P����IL^��>�'c5զ�tތ/Ɠ�w�g�rU�Z��1���\�o���o�IV�w}ɼ��A�3<U˙�K�o�X��b��`-ΡDˠ��^�,{]\�<p'���\XFR���-S\�2����
Zǝ>^�4�$�bg��������@�%
��E�P�~L�R��@gJȰ���aB�l�!�w[��L�-a��3�Y�2��o���1AF5��E3�zq�H��5�+��Ԕ<�D����,��U��T1��|�E�:B�0V8��v�9*�%֐��?�,��1�Od�}�I� vtj����#��m�~1#�� x� {U��vK��i��	�H�i�$���L����Ԥ�Rl�A���8�#�B]�qBc{��]9Ư�7�{�,Ս���o1xA{_j�#������n\%p���u�$HYd3#���Oq��.�QZ���G7qX_�D�+���gz5 ��I������7�W�.��ЧK;�AdX�T`��<��{x�)L�* �9����H�ԫi]�U�ص%��C8���9KE �~F9"8H��]V�p��6��1�[�r<�0d�W��u_�z+�Śs"!W
&ۿ�.ſND���V�ɰ�~T��#������5�(� ��g�s`��� �-Z�&��B��ځSM��tF&E�ֵ�xt�>*�,�Lz�D�60�����I��.޻|h]b�'���"ֳ��h�1�����n��ʻZ���_�P#(���ԩ�(eV�9XD��O=�H)y`Q0ݿP����`��fٟ���/��U�d9ØF0����4��q�~X0��F+ҸP��xp1l�خ�v�:�{ٱ�}�8����l:F���"3g <}�ZJ���?4hr�\���@����o�uM��5���Ŋ�!���v"���G=�_F\5�5�b<�F�f��p!�C➄G�c�4.Ni�N�D��p���1U�AF�[w� ;���Sl
h�������0�I��7m^� �5)�EK�粖�AZ�R�_|2fo�l���s��@|���,0��{%�N��:�#�!��lĥE5v��r�Id��H�h�6�S��?��6�o�"��w[�����4fJk���*���bp�iaJ�Bf�6�6.�5�Ҵ?�i3��r�m���Y�&��dVR�Q1�e�k��T�<�

�z`%�X��
|�60�p��P5�/j��E���{)��oe�e5���И-���婃�bd�'9c��S�H�yNX yw�"k�t%���x�(�t�T�i���P ''L��i�����Kk�i�'��J��
������bU�\�H�D@J(B!��#l�KPҶ�f���DYij<��w�̲�J�p�A��_	�s�g+o��dS���H�$1mزz�GY��%�Z׃)�ƌ�Y�ؗ칼h�A&���h����E���:�ip:���#�Z�4jQ�k�]
��%��q�.����^��n~a��mh��?�C/��
N�u�V��aG`�|�Ŀ��+n�i�O��xXr��]VN�gm��7�r��56/���OR��|*<Z�[���qfͷ����b����k�l�D�U}3���]��f��i�ˎ���(�9յe3יC7hq�,�@�}��mc�R$�Td��k��{�+r�l��cz�ݬ����{_�R$��U�]�s)e�;aJ��J{����*IE���n>(�US���+�	��n%��r���>5`��2v�2t������-���P��md1�oT��:@Ǳ!�"%������B,�F�:^.A5�E�ˣ��R
a�z`1���d5��O��
�6|�~4&H%���@蚦�[�	��GJH�գ6���o4��=i�詥��N��Z����o��-����4�c{��@$�u*ޅ���u$X�������vE��Ybe���^�e)��Tx����jr-n��<��/k	y9	g�_�h�:��pzm���ˆ�w>�&�I�W���%5u|�N�9�խ���x�,�Ӏ�����Bj�}��Ϣd�89�D|�s���"~Ad��uH����!������S`�EJaa��O���>�8��u_��"R��;qAEf����9+��nFQ�&<-S�(���<�P�y����A�廈� SR+{k��ȑ�9�>x��b����	i������ ��S���j z�O�x�E�n!���S:��w�޿yb_�l-�K
~�F��I`�w4�N�>�H�n[5�B��yF<+B�Ջ ���n֘��Ɣ�gY�*�UQ(�:w����jwPͭ?� ��D�.j���?�l.��'�e8�S��8ޤ�8LXNq�D��;4h���E~��E>R^�=A�ՙJ)��B@� �߰���?�۾��S顗���ǹү�L۪AS� Ⱦ��W�;�S��!M�mK��V?�\��P
��yi�ɛ���\�3�A�h��4��⚁1 �۷��b�~��� �i���R*�;�U��BV�L ���D�����T8����v���$�&ؚx,qDeZXLW��(��";�~�Wk2��T��1j^r��
S:�b�2���֒aJ�eN���JEq@/�]���dB���=�G�$�&"�.���JPx^{����qJq�h�=(��Qּ䩯'����������K����"I�C�L(DX[�mX���R�������.?��_��Gp Py�=��Z��������{�k�w�/�k�E"��o�UP(�L��<��H��4�p�!�E��0�>���0�<p�����/�E��o�W~��*���D��$ȵ=Wr�?�RQU#uBQ|8-�/�8Ŧ���^�t$^�@|pw��X�`��ayfzo%��mE�0Q�2ρL��f�B��f<`:�EY�|nHO�<cɸ7�z�Ps��+�������=������w��O<���ٝi[��k������A7�k���YJ��Əvrf��LC�&�N�TCS�����C�8^_ꨱ>��:��z������m��N��E�@\̟ˤn�k}����6���d(�b�{����Vo_��l�j��5�f�7٧<�k���M�:]��RjO�m�B7_ztB��~��dB7_2bϮ#>��1QeSFX�+��l?P��U���X� ��y���� ��]����+��LZ�c Y���"_�)*}�BB��|ő��6p�-/��S�
�E�����ʾ�?G��5��V��=��>%�~<	3�>W�GT�ޘ�$W��d	;�}���U�q�LiW��`�ѧ�%�R�@d����"'9q/�pZeFDP��TO�e�*D̫r���Sų���k�|'G,���ݰ��X���*s"��c��,h6�x*�9�VOx12ZYq�4'7�*�]&� I��c2�H��I���'��:hsl�y��� �������~��E:;T*�S=��Xtm�)<�����^���m-��V�_��"ب���*?��RG�n�s�����W?�"A1o��(#�h)�(N)P�؟q@ı�1��4�>�6B��8偝Cv��p	n���B�}ȴ�`��H0��W3�=��8���~���?6/�Uʇ��ڣ�NK!O�%�:re��(~�Ɯ�&����TW;��,������O�lG� !2h�z`�T@=���e�e��n�^���G]>��0A���'�{ϝF5��K!�s-��ޟٷ��6uxz���N�w�E�!�:�>�a]����(N�8;r�l��:�@��U�+�����MH辖�aپ��,�Ѿ������h� ����gt7��c��Ņ�Q?J�8?��X�p!;<��_���ڪ})���]�X��^�l��ZtX�~1��	�H�X"�sg,��@�\,s�w�����:�Rc@p|;mƏk];2�����rF�8|Q��ܽw�È���4�Z�K?Tǁ*}�yG�W��}Oz  B���$�qJ+��C>UA����c�M�H� h�P߆�e���i
�N�;�T͉��s���c���As���3W��Y�4��
���3?gZLh_�3O}��-Zg���ѐ��6�E����;f�Cn��GX� ����L=I&p���|k���Q�3�wsqUt�� ��k<�I_{�$ѐU|`$nF���V�ne�����!���y�#��c�,R��Q��{x_O:h�vTA�JR�9�REw�t͆����wt�o"EC����r�Ǔ_����T[Q]W&d�}v�x���SqN��n��F}�8$�Ճ���w��L��@k%��X����G�)��.�J��	��֐�ã�@ʿ,P�,Qy�QQ4Š�>��I��xO����������J�?燡�����o��	�_ey�}��*�k��R���2PK��|#�D`;O���O��G�X#�[
�˟��Ua�Z�m|.+�I�z�����W���?f��7�ǀq��h|9���v���#Y����K`�p>9���e����c=7G�'�l:��ݴ]L��ݶ�ĭ��.� ���D_nO1=�{�5�nH8G��l��L7��e��m+��=q|��O�t� z�u����mc�N r,���(���_�@�d�?|ٺd�Y��#�.�N�I-��q�P�#Ӽ����;{Ʃz��6��u%uercXoO�S�#,�� ����!�9Io�?��W����>�W��u� swʑ
���~�zCuP=0�֔wc9[�X�Z�H1�Yw��ۆ��!��ܢl�4��^�ܦ���Z�ҖL&��̂e�� �:�z��Z&���Z�RF�C�߬>����u����m�ꁪ��~�5�s}}�8�HY�_X�����hDj���uZ��� ���ʄ?�I�asmV�� .m��W�T��@vBdu$��үj�rJYΆm�������� ��:��'��g�ɲ��b�g��lf����t���
85��=���!�^�����(��p �ݔ���D,z @g]Y!T4��p�d���P�N��4�b�Ut�������|�Ȑ�2��(�z&TZp'a��7G��̥���	��T��D�G��zb���y��Cw�I��ҮI���rx������8�i
�m����|S�����lv-�1�1�pF:q��1k�RB[�(�l��P!7s>�L�S�-jRwN���Qo�5t�=\7i�iU���Per�L�g��Ov�٨�b`������>�}S��Q���Ȣ���{��Ti�$�j:�N�5wAv�cM|BNIu�WF76�jt��k��)Q��E ��?)�J#zq2sT6[){:z�թ����w3X�2(�����/S���Q�a���1���v�HL�����I��J��	d����Q�K������tqx3�[���rn0�2��v���&��vf���y�ˏ@-��D�-ʸ�/��������4=I9C�	�~&�}7�w8K�Z�#�Ïh�Z�׃9y�
Y�$h5����Ҹ��Մ�!o{ԍ�����o�[.�pȣ 3�"�6\�-i�hZ>�RE��.L�������>�v}t��SD^����`��}�j�(�Gs�?D���������OxR=�?Y�d&m�,��[��fBv�E�f/���	���rF�?2����ɪ��хV�5���H��U�PgiK�����,ٗ��};:�MK�B�L��� Z"�d��z(y�+g�ZY�eW�I�]��=Ч'�����o���`x�������*����u�>�ϯ%�خ��Y���Yo���L ʣPy����"E�	�JY��6� �`X����B�����\�W�Fv�B�.��p�o��sC!����|9�U(	��@䌻��)�X���~P�<�������8����(�I6��5��p��3�7���eч�N\ߌy+ ���)�x�b�.�VQ~o�~�q�N�r_�KM�<8�-�!�i]sI;�ܟk��q�]��E�t��-ݩ�;���%�M����5��H�Ǜ��]>�h{H0�$�2���x�=���A{^�U��х��D@vK��Qq8�h���!Y����N��9�V�3�uӎMK��H:\���b�]��??@�'�m���d�)޹ i~q$?W+��?�8���?�_��O�S(�ݠ��S> �9��H�Z���lAƝ�e�ZR_�]�.n�:܀�H�jMv���̀5'hU�w�
QY��$��9A/CtPf�JL�<��!��f��L~�5�
�F͚u��3y�F������&����̗^ i�n����?7��,��z��%����|>�p��E���k�#w1��ޮ��A	�����-�`<������b��>�l�[���&�����������'c�=x������]�÷}S���i�U�־%�k.�54�@����/��J��/��eR�M�Né�}Ń�|4�g�ڟ*Z��N����d�u�u�:b5��L�y^sXr��̿�|G�ϊŇ��ߺ&M��_rӛ�l$�	���)�2-��������$��.@�Oץx��r7��ղ�KL^@�q����Y����G�)U?�Wa7�=����j�/~cK�u���B�����<��i)E���%Ưc<�A.*��'_-���F�s��%c _c�r�>>��1��z:��+"�N-+�ƽ�s�f�|Bl��"�ꀎ�'����߶�X�����R�o��nb��~�Q�3�y������ ch>m�M�^v���$���E��Sa^\v%Ж��rL\�؃
�O�C���^b@�1څ�6�E?���z�wvq�f��,bq�ݧC�ƞ��X?`m��p!Z^�Mp�M�*�!�H|f�M�iU@q�����@���5��!����=;v�k��}�o��t�u��P'�O+k�2��f�c�i��Y��
⬺�����������}����q�nr�x�������ϖ�pR�`��xE���\���;V)4uA0��!�����m�.����OE��H�pe��wE�wh�W����L����Y�h9�}i�tjD�*$����3���U�#([��;�a(���-2L<�b(�b�P�7�?  �9��5Ɯ;��\����JR�g���]K�P	�Q-Aĸ8*P�������v�;�~S�~_!%i\�KZ�{��u��k�b-�3�۷[��\Q�I�7.oB����Q��Bgy�d�].���]�qt �ɑ�MOy�#=d;&#��߻��/̌|*1ہ�H�r�h!�ݖ(�M�� ҄rFM~��e^��O�P��E�@c�'����µp[>��_z����_��FQ	5_/��@��h�S�<X�G<��U:���?~�� �"�ȓ3�j@�7%z]@�0�^����53��U-n�D��'G(�L��>�oO�
7��y�J��ئ�r��a�CMK���'8���Ht�W
��_4<p�4�[�K�(g�˔c�e��`�F3(l�CɆ��d�x}�ڹ�.+6cͿE�6�=6���jeQ�i&`��1�g�t�<?%�aj"����W6$#��\_�MH>Ĵ]�V�^9��=d�|��#�Нu5�g�X�?��GdU��r �u�,+�e���.��+��y�q:2_4A/�z�	y�Kp"9Vl�� :ʥ΁���$�N&�V�'�@��Ƭ&a5�C����t�.�2t��zn+/���F�F�X>��: =��f��͢z��y�`���#)��
@M:?��7�?��㿺_��Z��P�aD�@4Ot�v⁁�	�S��R����2@���QX������c�<���%�p�|����\	��a�,Es����:�{^����t��n���"7�*���&��d��m �7s+�&�_�5<̘��X�K�J��~�>�bFmɪ�'���%Ӱ\k�"a p�@b%�C�.U�(&�G�G��?5�&'��F�Q���YB�4��ݾ�����3��^�O�4-�A;JD���_f��ٙf��0
�2L������Ĕ�M
p#�~H�?$��)�@��k���܀_��ڋ�,RNQ�(������Phbsu����L�|�m��f����鹦Eʊ�������6wgph�ʈe�Ũ�[s�dS��^&�7�d�������A^ �G�鉅�:F�J}�F:Q�$�ac�%b=6��EȖ�:����eA�)H9+��ūI��i�Xv}���`���
$ߎ�z���Pii`V|�%i�]�v4(6#���M��6񿕣�V1u֗E!-�E�>JVǛ��Y6�ymM"��N�*�ds�5����i�~��p��&v-�
��3H���B����a?:~�մ�19�@�����qX�i��#�K�5TF�a��D*����M��	�ҿ������r�<�CC`�p��RE1y�Í�[�͋C�B䕍�KO����'�HJ˭�ԮS܇����2�K��1���{�n�����A��ij<|�ύF��eg��e�F�h��ٯ����5�Jy�Lx�7i���}���p��_�̳(�&ND^�Q�V��r�:W`8h:�h���%�����{lH+Bi�s1�Z�^����q �(��t�Ԁ���@��v�g�Y�s DW�I�?&'ܻ���D��>D
� �����^y�C=�,� vAT���-⅀��~�� ��;��<!�ę�p`���k4yG�hI��&��vg�Q؛����$���RE.�����zx����m�ۛ/��%<!19��{S���%�a�̛����N��-i�^��fc�:x�b�3{�����k6�bmi~�tZܑ��()�Еg5q�HXOZ�q����������#�z�Ԧד	�l���w�"�#�]v=��'�O�8�X��	�QҴ�i�(�DG��`s��͑-K�y��v3x2���d��8c7FY�/^��?%GZ�1`�����k�-3����!�u��F=|�D��].�_ҹ�.D�
�U��̓�� `�tZ�vq��A�qOL�\dL�??tS9٤�E'ctò.6���	�鵦)QE,k��O�h(������*�x�?h�9�u�U��>������K��a0���g�߈�g�S��1T��6Ҭ���`0R{�����yT�M���~�p���o���ϙ!}����v�@�'J$�}�B/7��� _t�U{�{CS���R�{���P��Z n���W㯘����?挵|�4���9����5���+�������u�Rޤd�TE2��/>��t���t�
ԃ���3�u�A5��+��7�����������Z��*�ur#���V�!�D�Ijh��GK�F�h���l��^B(Js%5Ԋ<A�fXVC��o��MR�J�^�LFK��77ز��v��� �Tc!z �ҩAU�s������8�[���H������-.��V*�ʽ.R��J>�[�̺�V��;����C!�'�Ac.3�F�q�oj��<~W�W/W%���m� �G�L�9�8��5.gh��y�ke���i$ڴs�p{�$h��S|����&�ČB~>�թz�{7����<��T56]�jKAx��7��t�-�:��1b��U����"Y��(�B��u����f_�C�\�ik���4A�)��v����4�����º����ͳR#IRȖK���ͧx�^Ey�709��M2hGങn:��B�<9Bg��lG�e����:�@z���J�X{�? J�*��� 	�9�0lb������~3:L�d��VK�eql�&r��.�H����,[<n�9o��5<ɃG�\I���
�9�0�{n\���{mP�x��"��h>-������Tr�T���ҕ�+���Fok)����L�n.�sw�pZa6��T�#"�D�a�3����+6�O��R9��g����8�4�T���KxͮMU��{T�y�O��4��0����&#�g<����?�z��;�l!1��&�Υvñ��=q3M�%���FN�Ă�;�rx ���a;��Փ�F�|��˜�}����_D��!}p/�����Z����򜟦\m�eZ�E��M�U�R�%�W,�춒�ҦvT�7�|@�{�J.V�Yh��&mK�oQZ6�{N �K�wļpn6��N���F�<��-/*Y�>�țU�z��B˖��H��1��ՂB��Cw�Ա� ��o�+��mT!G�������<����r���hۙD�� u�@��J#�uMi@�#g��= �����_��n�j�pI�w���K ��i��zNjGo����ap��%�rb�龺>w7a�zYl`Hl��{���`����7V2�܏�,˦�G-Ke�[4n���\���䌷�A�Ř�Yf M�v<�.%B�ߖz�x���lh���Pp��UJ�p�x�Y��&�C���ʃ��W�7k�֋���5����z�L���t�y_�Cj�W�`g�9��
tI_1P���������h:��<���J5�72=��I�iD#�❪�_z���3�3>��^�p����0^��+��g�\H�Cg��jx��Bn��J#��7$�_�lzJj�g+�2_�-Ne1_]??��+:S�a6Y`)P;����;6�;���݉�*'���~���"���Pl�d�Hz��=�b���il�������h,,�z��ת.1�A����s�*l<�]����6�u`�x��D�4Śi������u�L�!����c���`ĵ@�ʼ�7�B�!��R�P���uq'�"�M�$��� �6���)9b�<�N8�Y��HQ¯8�AE>G�%���K���iL���D;�c�Cq`���t����krv�W������jɽcNUvs�6�iE�#�t�PA�O��ud���!ZY��L��%~����\꿑x�t+zW�Ì0����Hգ�i雬ǐ���Y�����m�Q�7�O�o�ˢ�;�7�Ҫ��|Z�2$FUrp=o����Of�W�^����0&�I{�^@A�#Fz'��0�q/!�K���:5���z:~��p5�ra30���A���=^:L�1�������s�q@م���*g8��~Y�E�1��+�ߏ���Ak�-)4��6��{8Q�����M��>�3��	V��!��L�Yf)��$��V�DT �)FȔ� 2�����I\)��a�xP[*�ws5d�Of��yp/��=��o��jąE�W���a;g[IP�۱HAd�w���@M$���P(m|"�.)H?00j�F��f)�+'�W7�_g6fɩ�;͜�:��L
t��x��ͬ �&A%�B�$iq* k:�B��N[2�K�:Gn��<�s�r�o9� �����ܙ/]lE����94W�)�)T��E��;��'p���
L�-2E��E6�#ef�z�^��@֎�9,�A��)>v��n�&OX��R�e�N|3$@��0��ݫ��j��d�O`�;Hq4����}U7X��^�B�D��gvؖ��2S�%+�u�B�H�c} ��𮉎v#W����~0�A��9�[��-%R.�kgMX
e�(cELh�x�b����D2c���.�����I�T6��eSX ��9���h#��(�J��Wi��;�����D8f�<�~��!�\��?�[�A9H��A���W&��##R�}gbIkH�"�v+�Ua�������zCDsc8P�}�)B%�1�[�{pz���J`��:�s�_�G
sp@^m�2=�=�U \Ϯ5ଐü������"��I&F,(jF�A��_72$)�xS+�)����f�*��o݃RJO��4�г~@{��4xgܭ����q�����3�>2$�dZ&[DC_ƶ��
�I���z�nFn������Y��Bk���)��܏�����Gc���+Y2݉�� ��� ���dǔ�ȅ�9�ͭ�c�P�}��;>#YՎ�U������Ѱ]=�0�e�Y�K�+�b'�ζoVƹ u4��1�R��-��p0;�%��Dl#����:��1�?�%'�%�"ؗ�K��ʚu�Lq+�2,J3�'�1�B���Z��H����I�?#4�Uh����5����3nka���:�,�����;�Q���O��<�F6_x�Z�r��%#/�!#|JP{:�l�[朽eF7�#�QT*�[�a�|1��S��5�_l�2�(.\�V5�u���.�i�TP��5N�T��C	5����ㅕ��.C�<�b fPV��[�Y�{|��18��ol��!	����i�����z����}=��M�Fꛌ�|�^��fn��J%�ߑKOj'ys���PnMh����R#ڀX�1��-A�(�t���u+�/Z�̡��`�Y�Ky���qyd�Ci ��!��ctV�i����X(�oͿ�;�tJ�x��A��bjK����$1��V��x�qR��=!�
g1��AiQDP2���2w~J㶐q"P��V��%�=�n{|m�Ld�b��"<e���
���&�#�U�o2��6�U�`�e	y�37�~T����һw��o�]�IgԌ;�l/�Ҽ�w*�D-��n7R�צ�W�@� d�26���Ʈ���X< ����p��*���s�E`휘�9=��l��zc\�, w~V ��שS���7~� ~q�R�|�*�y;be�XA�⌡��������q_��������v�K%B�n_o��a]��\<�O5�C#��/yI.i��a��ɑ���:�\+�ZU���#5p�>��}�D�:*���㾯g��X�_�~i"�_!�i[��OIЕ���j6'g�?��o��WY+ނm�Ǳ�����1-O'�%����,���q]�n���f��x���)���{��?=~�4���s��㲘���F��a�e��5�Kmd/7�����.�|i[i�i���I"�(jb��y�Ҫ��-(��ڢ��=x\4�	��n����g���鿦����/4�k<�ue��Q�
���5f�.gͲ%į-�uy
��歷z�em*H��|����w�T�/▨�BV�+	��s���meZJoC���R�Ү@�ߔ�@t�*���w������q���}�|�PѕU}2��mE7�C�&�Wd�֔���OB�<�$�2�x��	��f&o�4���=x	)M�51ZjCx��2��k��r���l�
��t�X*���n/�9��އ�+�+�0RHAȴ�|	>S'r"���r?=���J�w+R�WDf�fȞS�)�� JD��\*����/��?�&����'�6������%uj$Y��b�k�Uح�0��������0T���8�b����WC�N@��X�J�GH�������r�ҷ��BJ<"�Y6��	�h,e��t��A�,g��8��8���B:�̮ AQ5��G	��iܕl���%a����fη/�A�Û���0�c��]��]?�s�p1H���P� �q7ML�uu'�*����~rL��(���3��zc��X���|���e�i�Q��#�zM����^�eNQ$q*�M�|� ��hc ߺz@��N�[^�G5��.�9�dM���<BF/�q��D6��h��BT
\Ї� nr}?H�G����`}�B9s���y�(gG��ei^v]���iR�N@����)�8��m"��6:�(�t���J�ʩ����d�	ijи�h*ɡ%�M�R��I�x�)� 	}�#�wX�pv�G!�C�isR�(g��'q�t���f�\�����j�vQ5����AN�*.[]�^���/�v�=�&A���A��q9���5�:����ٌ��+���4M![}����_�S�E���9���a�~�0�� Q�~�.M ��%y$5TG
�*��u�2,k҈��l�_5����ח��l^)��t۪f��L��_גE�U�Z�Qc����u����8������|)���>M'��\�@_�|�ݒk{2�%��E�-ϝP�Xx.FÐ��Z��M�I0����=��k �p�'�|�j8V�~�s���n�	����� \1#�R���?6�&�7����aX�C�EO�P������9���v�� ��4w��\���zD �R�"��3� �Q����.�T�Ԇ�g11�fel���cSi�gs���đk��R8W!�ͅ���t-:�b�ܑK/v��w���ܐ���GV�z�6Y��{�+]�n�3�(�3��')9vD��`�����x
R�Ya&��_�ddۼ��J�!j>�ha�˔h&��$L�g�q!%m1���[���������W<�/����w�����~�k6ڬxSxz֗���XŖX\��E1Z(�a�����S���X�����|�7t4y������=��F�R,�F;���ҒpYgz�!ޜUb�&�d�@���V؄ ��>ܤ�[�����göR���ŀ3��S�ڈ7]<Y�sю���\�r����Bd���۱t����N��et��Sh���L�(��W�Z����l2��I}��F��b?ѭ��<1�'N< 	^9@�{���(א�������#�Ͷ8���Q�C1$� �A��ºu7$n��?�ʨ~4������%��gӕ�QK�A^-�\�?�m��t�>���a�@
0@���?!~��Q�5=Nl�]�"/�����"e t�>0�!Y=�Vr���������n*V�Z�8�}�ǣ�q���b�Wpn��w���W�0؉���m���|��{����I�n*P[�Xtx���ݕ�k��n�����9�[= 
$�cO�⓺��q6���#�|̆g�f1�X��84Zx^���ʤO��Z΄͎J������C}�u�?�>��n�;��B�F9�@�L'��o�]�$=�hݺ�D��'�@��Q�uX �v�Z�:�Idhou�Vo��!�ą#[�_��?��]j:K�O�N>��D@~��(j;�U�B��4K���#�ԩl�SE6�:�T�n��?��Z�e@��R ZW/����vz"]���n���2(^��̓_#4�R$[Oָ���o��~�ATi�x�da'K�}=ȷ"����b�3�k�&��V�t��N[�{��,�$ |����ĝ������~ ca���׷��Î& p�쏒�>�ʀVg!cI��r'�l�4���6<��yG�
������\�j��-�c�w7`ALnO#�I��mH�u���4th�y٫J�)��K���.�����[�`u9��,��4��ݰ��\�<���B`rh9.%|pm����h����L|J��b�,�Ɗ�@w������^�*���s�Uÿ���,4�o���[g���Vd�L�N}�^��:'Ne�c�<t�l�^�B}uD�d�����1������D�wM�wk!�9��'W'�*��6�d�d��(����{ٲo�`�&O��yX�O��������}U4��I)w�V����� �S�\�����z!�|��{������Lj��p��y��#�O8ۯV���Z�f�EB���?hG�f�o��+`G� S�UB�x�����R"�O�9h+U�Ig�r\d��x�N���/�G{�1�R/���Izg����� �xi�,�u�B��D_���c����M#m����g{�t;��f�����rE�v���Ž�F�8�"v-%z'�;Yoب��J�Pk��%�cĝ����s� u\��y>���޷�ц�쓭�_�1�՗ᣰq|���Y��R�� �Pw�!��~H�;�e���Ԝ�/$�T�����lݺI̺�Z�Jp4p{� Γ�'$Cʃ$N4=�t#��5}?���Fp�9�ښ����f�(ۆ\�;"����s[>�����N�:�V�
<��4j���/�?�gS0�/����wwU�-2N�2F�@��X$�Q.��6-�>�80C���mC�UI'�`WO�H�i�;�?'qF�5ѳJᕁsM���Ő1���N���Ŝ�0;(�1�r�g1Ib�T�7ߴq~��B�P�ݕ��(��P5�����q��������>�qo^{�Z�C����~����>撆��]ȏ�v�����+�N�vv�p��u����gC�]ʹN�9�\��ظ�f�����Ǝe��v�t�.=�ռM��(����Q����%I�Y5ER�Q&��]W��we�d�[���z�'�4����T!d�b���+��@�ѥ��h|���jk�thⒾ�v��*j�@���7E���n#0 ��G~�xG<�`\Y���}v���nD������K�	���4v��ϯ������p��ٶ�˔~_}��4%�W���,��Z��,ƤJkaH����.�:�f����L&>I��³�Q���"{I�9���ps�@�y^ا!ٿ�֚�R�,�=!f$�>0x]h^XMtۼc+̈��n����:]M�2do����T�9[�ر�����*�g�k/���ރ��EP�U���,]��G�͐���xF*�%IW<X;�� 3��bPW�|�y�������k�1�߄b�@������iIt�k�9WM���PL�E��j�*$@�Ղ�ღ�~�̢�l���%�����-�3�
���^͆�T��T�ѥ��JV:%�;~^	�f��:��̍e�e�g=dol$mF�����9X�U��Lk�,8��hi#C�#�oP5%�$I������a��G��KR�������n�N�����}_�y<��=��Y���W�U@�cHy"�l�c��|^6"��#-��t?7�䱄��4Nt��.��x��Q0��0a�a%�{UT�_@P��E���*��ג%8�g�&\�+�喳ԝ_�4:��S�o�b���Y���(I����bmN��|�B��\� �j[KT�!롯�6��@��%��[�D�z���[��4������Z.����𳤕�%Bϖ�����B;��Դ���G���!��vP�(�P[�ج��_o��u���s��&��k ���d��D.E�>fa��8�X%,]c��s�E��!`�㌧���g�U��h�3��k��)��&fg�4��H��� �R�kCX�%�sA�%��u!3������F*R�\x[[�ndC�d���â=���b����c�!��}����ZB�<��O�|mQC솧�}ZC���F���K졶�4�Or9I��6�p��ONWX�n4��"¹�D=�P��+��X2B	�3�J{}�y���pt��'r͚"�_�`)XR�|��;���KzvVS�7fi��AZ���������Ө��E��z�8���=/��\�?IOgrq��@���rgj���l�f8v�u8���[;fF4t>���BQB�&�5���W��I�m�v�ħ�m�K0��/.'G.��}
��&����B�W&`��?ʟ�A�"�瘌��@�"L�V�6t����GSLD�sȋH#���Y�1\0e���(����gJˁ���+5�����k����wG�i䇃@�X9��O� b�M2¨�&�%�B��yU��z�)�E#�bOX��` �p[�*�H�;-����eڤ��T!���?>#�`�� �}�Fx; ���U�� Y!ƙM�_�Ձ~�1����-5�:,����l)����w��
S��,1�z���2=��a�!Y�Ǘ1�PAx�]�$��?���|����O�ڲ
w��$v5�p8XY�>&��&���oa��k���洰!z�4��$
yh��E�Z�?���!��C�]x3SZ�e^t��3��6��kb%��]����a�O�cm(��omľ�?����7�y��� ��4,JԢD��m�]��$5�5LƉ�Ȥ"ػ~�Z
Iש�`w�u՛�w}_㙃��2��eO�u� x�$s�~�h�6fs�:ͺ����h/�b�%	��2�d�Ō�(�'�/Ǖ�~��;08���![�jl�WA!w,�ՕIV,��Fͨ(WwoO;�QI[�'�^��7�����C`�Q����B�F����m	�OZT=�[Ƹ��}��-jyRwf "m�`%dLjȮ���%��dV�7r�g�/�46��'!O����#�%�8�y�:B���&�Q�$�O ܁�[lKũ[;x�7��D����`ƿ�g�@<�Q� >�
�;dpK�谨�
m��h��;!���F�f�6�)�o�������k�D���a�w؇�X��+--���'7����[I�~_[8 =��n�h�*_`
U�Q��p��N��S}���?F/�~Qc�M[oN��ŬZ!�v�Kg�}�<v3���x ���%T{1���)6pA�O��Ok�W�`�՟�O�5Qdd��ZG^#,��A
3�Ƀh����=uߣ��1]�"dF�>��P����P����╙:�.Cn	�i۽	V�À���x�`pW�g���*��5��>� ݭϮlq��[����-�������;}�6�@�}���٥�Qx ^�[6�fOQ>m�4nP��j(@�cR���6�;m��)l�b���P(�G���,K,��)ܜ�q�M�����>+�e�"�稙�Y71f\"����B�����]0���kM�������Ҵ�k���Ǝ�ʃ����1\7	j�x�G��ʬȋn�Ȑ��WQH�b����Zh*���1H��&Z�q�_/Og���y�p_�����l]+p�[��!zwV��%XLnjY��=6���������f��y�%�PR�=_k�/��|>��sA˒�)5��o.�R��l��1�}��� �Y~HX���X�+�Tk���.�a�)F�PyM~��e�v�:�F����5����>Mк�,�̆���݇��h������{�3V�����ZBT"d�Ɩx)L��k	T 9��p�lA�����U��C���tD.�V1q���~[�>a��h�DKN���#�Z��8%M�}�w���6�&�3����n[��f�=�w�'��������q���C�;wNƾ���>r���O���<ٳ`T��I�
�<��EP��rbZj�g�?Fmлm�.��?E��o,�D1�q���~��;i���
7�j0�����O�N�8v-�%�<� 6`�~��W��g��hGU*N/��V�F,K'ʹ/��}���iȚ�qW���ey�DX&hj��.�w.S��qb��	Ƌ��:_���]�9�r``�#�zmA�(�@�.߉%��w7�����������2a�̽�s!_�`0�&T�)�U:�ӈ>~_��
Հ)g��8��5#fF'
�����Y���q�J��ǅ=q9�����4pO���P]uH�^1�6p��yW�.I�iڈ���L�d�#X�1�����?�e�.�\���3�S��;$׉�Ν��N�YV;�K(�זܦ�������t6�E�'���E���K���R,^X�����_K�zo8���������IQ��(���$��v+V��SfM�q��w1����|Q͞�?,�%�C�/��B�5A��tG����
��F�`������x�,)
�h��<�|�-���o���S�����&�W� Z7G_�4��hr���DM�W�^H=b��wտ�G�r�1��En�Shc#�]9s���'�:t^�*Xh�1y�z=�fy ���#ħ��R�8=�pe�i9iY+���K%� �ʦ��Q�f�m�G{�<�}�{��϶�P�WWr���T0�Hܞ�}�keO-L[�>Kbݔ=2f�^o�~6t|��>l^�Kc)��˂"���W
@]�QZ�a�,���?�.��0�$���"�w�;���+JEl�����(��C݅qNIδ#�1>�KpCzG��C�|OQy���S��f���N0&�ʡ�V���2V�:꧗�}�zT�U��N='�^&�"X����Շ���L\ V�Q��jօq���w�#Ƀ`���Z���:e����?_���/"~�X�JX:�<w�fhZ�����X�vB�v}Uf��$�v���B25���Gח��/��o�N^�+)�6�h�'4׶�fP)�Q���u$��N?߸UG�����0�Ί�#b'o����������A9Z�Rd(�p��0���-Rt������$:��h���&N�)�$"�*:��0��Is���8T��v_��{�����l��v����$�[��m�Ƨ����{I�*"!��1ia��F/���ow��xH���wF�od�l��#�����R��З�v 	�n�pË��)�ۆ��j�y	��ni�������*F�0����j@��sΣ�~�4�5J�li��J���#�kĀz:�O�����G�ӫ�h�nۛ�����/A6$�B}tEY빯�j��%��-3�&����Idh�*x��%����RJki lH���su�Z���Uv�]���Yg�5��ξC��-/Sѹ���B5HXO2.L�� 9��7ɨ��HNu�V^oK�8�n����r�����G�9�dr��nhߪKSɚBA�)�u��k���.����NfVuM:�-` �x}��yz�C
	B���M5ut�� �Io�6�?S ?���8fo �y }H&�%��^�3Z�w�eE����t��������t��lk����Y���0&�W$�)���&�#�^մ���)qW���i�յ���������T�����mE>�� �	V
J�˫�j�sR��WM���5������j��;��X��ѯ~��c&�Eّl�j���Y��6<��_�k���/�S�D,�z�	� ����֫k����g��u#����U�p˦��l���Z�?J���ʋ��^�(�@�[�-�Olw��$V��hy��T���пwcjLz��Ĳ�I��l G��*B��������`���b�!�W��ѹ9�m&xH��;NM�'���`(�K7�]��{�=�V�e�#�fE�D�����UV��o�$Lts�^�U0nQ��J���[����E�G��1�0%��)����R���n�I�sR��k���Y��\�Ɉ7}����U�3RʤW]Bs@QKb�+}�pʬ��ؔb�{�LؓO��
�P��ǅn��4��"Bf�
��,:Q�;�	��	�Q�B���E�?%� ���:�Ko>��v^ȭE9b4}��u��o8-wr�����o�M턼�⴯m�Y
���uZv����T?b�����ˉbA���0'oy��E�ڽ�|у^xq͓�
+�d���Mx�t���e3U� �ó��=������և��ɕh\R�X���ٸ��`���37��+F8�s`ja�����eB2`��cdF(���ML~�v�h+��E^S��B�^s�����n�o'8��Fr~�КA0��
 ��`.�v��� 3���X3�cc��X���%z���b5t4s#?��-i�"��sp�)���%��4��_j���]ͽ+$����U��k�]���@�gc<�2M��³���	��ڢBos���!��Ձ��ʩ���l���o�ū��`�^5���]:�u�9���m�ƌ��S���d�q�p�	��X���mV����r+�
���=~<}����"����0	��|���`�$14�d�y�\�1j,?����)�h���7�� �̭q(�{�-�����H��;�G(�wڷd�\� t�@�]���MEgr�Nk6�T��)�e?�f)�%S���j�Zȣ]LA�F}���t@z|�q����`sz��v�M�+�JAJ���3�ǩ)�d���9u~��9���Q��ܒwٙߵѦ�0�2���E_��|�-[�HߌYC���@A�W�,?R��C��`
����s��wnh�����}B権h�:(��N���ʆ`������V�n�ӞYh���Ҭ�Jê2����0����r��^���V9�1[��*N.sV@�"���xf�wʵ�$�(�����+G��4��}���w2�S!p��5~9g	Z
R�ݤ'!�-Ǆ�X��!6��1e˵�s�Ub��F!N{�g~-�-n��&_R\�͈1j�<t)]=�w���_f9�Zi�Q!IEu.�c��<e_���{E�Ɋ�7���Ǚ�PF�D�W}��'(�9A^N�,�k{�8�>��X�״�5�m�ȶ�\[��8�&��m��Δ��E��η�v�H�9Y���7�cY4K�w.V�aw7��ƄЪL��b1ұ�=~
*��k׭�����#A����&��CG�jGs�I����څ_|�-�;Ϋ��j��>���#�S���yHr��uW8ܦ6E�a!'iO�ufS��7�̺�S��3�Tw��92��ܒ$��v��x�i�\
!�k��w�imE����Li���]Q���'KY�춢*q�vf�Kⵇ8�7�R�~t4j<d%�1��z�� ��s[�/���3/������qS�A�7�0�/�YF��Ѳ��������2/O"����M�y��y��$�h-��0c�J�a�Id�v���M�j�jtٲ�.C��l�T�l����C�߈�hmm�eT�ELN]/�-U�x)�kC�)�Xb�ث�C{M:MI�5^��pn�5��N�!���e�X��P�t1�뵤��u�~�2�?���:D#�`ȳ6�%�=���Y�ƹ �#�WZI>x#�P9�&2	�=��ׅ��]�!2v���rS<���0	�7�D[���dF�@d#�+-fxE�M��`��SYD�v�'��Z9��uf_{�/.�Ts���K���
'�C&�RC�0J�1n�.xu�D�{4�����Q�	�{�����í�I	d�O:KZrNb��K��xݝuF����W�Q�W�'� �\����-�����vCbX�0?�jU3���9@V��$C��@s��>�K���]�u��J��w�d@�xt������T',�AO���n@�Z@{;��c��>�:z���Ð@�J�g�����Ȣ*x�v>^@3���j��T �=*�7{tla�Ȁ�Ȩ���1�p#�Ⳇx=���%�*�� 0�«�B=��e��2���`��Ee�E3y�T�4p4�;�C>�+�}{�Dn������B�hƎ3.��{ȝw�㚡֞CP�2��<��2/�ERƤ(1r�j�+ȼ�V�2����\0�P�Wحy�� FWIПU�dm_�r���C����	Vbh��j�L&�:<�rt�^���� ��Yxz�E�����_�.%�r`W�R|kX�?\jv]�ic��Ջ�}=�e��
���}(���yW�cg��B�=��Y�V?ȗ?�r3���W��V4�����7��YV���������t���#,2�ʚ-L������A���0�З�{�>
~9�u��8~� }�o�j����]��D��54�?���~��Xɬ���K{��fG^%�ѯ��NK?r����0(���B��܃�f�dPŪ'�~���_����a$���E�d�#�S�[��K�f(4^��똿&z���2i��`��t\·�~n����i/ލ�(����_��Z�5E~-&+/��뢨�������z����#��B��޼�[.���|}t�����i���b�x�I�4ga����u��$}~��m�'I��h��5r����4�A%�Z.�Zt�,<���t(����Ǫ��a��L8:e��!e��oփ�1�<`}�[>�ϊ������!��,Z�r���c���͜�1-�RP�����9\�-�WX�RE��壥PV�)k|>��/c��D:��CO��o��}��]�?&�������6o��L��-Ą>�v��:�|z�R����<�@��GW*;3�c��<���"5�Ʊh�c�;w:�{H�?H��,�V�]T����ŸZ\���7$6�V���*� (��p(W�|2cu�R���n��V�@ەa�Vk�|^��a��TM㿲%L�rn" /�Z���ܳ��q~>�!3�ULd��!ٕ]����J��Ã��)y�EKq�v���������y�3���$4�ȝɸt�"y[�͗�XauB�/�����f���J�����9�<�,��b] �.�攨��1ص?)��Q<�Ҳ�vO����Zw8C��Dt��}+vEP�kN�&aZ$i��0����Q=�����R H�7�ϣW+���I��t�N�	ϖ�r�,���yW������f
ЫЅ!�GJ�� �Ǉz|�\0���@d���2�x��~@d���H{8ԌI�%��������,<oǚ v���~��	6����,��'n��}�מ&���*���Q��jE�f�\~�L�y�F�B�;q��t�z�]X"���;0�/�VQ��O�K�pia�ώ�y}ڨ�{H͹���"�"�x�:|�|`Y�*���g�zK���m0�k5~jiri�\�A��r+�j�+�o !h$������#,��	�L�&���k�[ϊ@�\mOx��\���26x�q��c&K�Q�SS�sƙ����f��9I�.���hX��%gs��$�ѝ���J��ݜ��>�x�>	��x0Y��t�Spq���U��4��d�?�Qz�:)T�~1q��6￝�>�d��{DB�۸���_Q�!<����?���i�o��]�E&��W�o�>��L8�8%Rŭq�wQ�2�{ �g�|cn~�dBW�}���m�~q!���ĳ�\�'��9��R�Ul�i �gNu�lo� b@��h�BUi~t%�J�m�����#�	��p��j�x�H{������#�,�������6�Q��f���po6ڠ�;�t�"�(��wa��y"P|�M�GYфRr�|��h�6�\����ǝ<ä�{��ڕ�jZ���/.b�X{g�Ȥں���7����?s�<I��@�M����ԥ�]zg.!Zķ[� 6��b�X�Ǣh,/п���w��|�0�ÿj̭W�ed���1 GƇ|�NlYm@�,́gM�H�Z4+Y���,�֒���,�A�T�l@�V/�֯H� �L��\SM᳡����b����8��5 bCx����ɉ1;Ƈ�2�"_^�fW0K��c%"��r}f\z��B��S��)_�(,ջ���vҭ�'�k��y�lW�.
e�����R_4q�:	�cb���;�}�L��S�'rų�y'�o���z��^� ��~4��� ����C��B�c>�_ӄȳ���f+Z=�<HE0���1���,T.<�Zo$l��0�@�:�[�ضzAD�X�+��y����\�=H޴c)<I��\�^zq_Da�x�75ޢYd�?׍m
<ެĢ���R�A�Ĳt��s�cj�x��C$�8�����)��f��/>��x~���c�(��$�@���Q(I׍9$�{�`�ӯs����wU��NDz�cc�u5�FoWe�l�	0ߐ-�w�t�پp"1�lS�w� m)
oW��F�*��[c��� �x���Ҽ$�4۬xؤ4 �Q�s�w`��-���i_�g9���e�#>0*uL�=�9Y�p!�_Bm�`�΁d�rn΅�C�/���"fʏ�V��L��	� "������u������շ��E�+�:\$�#�]cp���)��k�6a�[���6�l�x����I��椅�c��2�z
�pgI�X�+H�Br$>#V�3Б��
˓���x�[d_�T�r��q���z!#O��Bx�� �Ua��2��V8f}��f*+4�Fb��L�HE��=A'ȝ���6����W�q;��h��J�dy�xqq���Y� ���lo��?�d2�~�p� c��pP��Y$A�X�	��B��+o�h�X�1l8��\�S~��ׁ"��_Hν�����'����k�c���e˻�IQ��V�F��$��얖�4_0����":8?I���|���@�po�.�?�,�C��FiF���(ib��!CӿRRk�[��&�=��o��(  wZ����W���X�#�ss=��];Aq#b}���ok!(�4p�ߑ�W>iEBL��}��n4����p����e�1ms#t*��"��)\��Q����[�C�:����|(E��%"t��?�wQr	��7�rT�d�a�F�� C����0�c-���-���I�h�
��{O<>��.m~�_'H�3���tQ���]�s&¬�\~UK� ���?��P�%U���řխ�@%'�K��f0>�rQ�!���O�6��q��>���uN�!QlH(I[)�uK��5�yi񟛓�uź��G�Q�69�2�缻�~���oVݿ�afժ���P%
���ce*��'����N�v+�T�~a.���O�O���'����we]0yOy�dJ3���4n�����	�;�$�1�d6����b E.�-�v���*�I��̚.e�>O�h\��s��> �.�l�tm)�S��(ᬢSO��H�~k��@���IG�����z���8c8'��]jP����$(��U�2�`6��h5��
�hH��3h�W	����X�d��7�����*���<;Ȓ����P"\�Q��|#�r���F��nK��� }G3>]^.��u�b+�G^f'�/�F{H�O$���_��߳�bL�2�n7��FTk���<w��7�p�}S��+<,�и(6�k+��av/hh]��a'���xVD�N.�R@�X,�OrN\p`cÉ8�@JC, 	�ZRPN+-HS�׀�������+�[���
a�s_�Rĝd<��ۮ'����$k�8:HKi���/���$��M|��a|��L�ʱ��pG���SZ��X�F�t��:9�)\��<�?xS?�@{��o���[5��%{i��r�=z�].Q��	�z�7'�S3-Vu�LQ����0Qξ��k@ox�����B�<9g~�ČҬx 5T�@p?����?$�*��;y��OyX�Ł�7˱L90ػ� ū��9<���Z%d� ]IF�Ơv�=�SXI7�O-�m��5��1���ᄊ`ah=bhni0��l�%%Eq��Eކi顴���8_���/{��ٱ��Mn2^��E�����r�P,N�W���n�nH���9K1�����Ҳ��z���8�������ѯ�zݯ�"Ib%N�Zً�����c��S6�,v�`������+z�^p� >�F[����Y[��E}���N���W��P�6���qv�4s��Dt*�)U�8�0���O�����w�1l�����T��:Ϲ�)j����>�
0�z�+s� zҗ}b+3��ƈ!�1x�3����8��)�5;�7-����r�{02�^�����@ۦ�(�ߗ�/�%�N��{��%��K<��9IpF�ȋ���&����U@��W�4�L@�o|#��V�yea�2�@�nkKo�q�'�-4�BRї2)��?���,v�2I�k9{��G?�Ja2�(7��!�n����*w�u�����u�[OJ���A��QT^��H�=l��ũo�"�'�Vְ$��������텒��$�=͋���ŧ���b��3��;?Y1�T� 1�f���� ���Y(���BO��`�O�u�W���9x��p#\啥���TK�*q�{L[����b�S�쒄�$�+�{�r�\ ���`���
���jsv����2���g`0�Y<1��0ȯ(V�A�ע�E̔�N��R��(�eKR4�er�%��$N���b���t��x�Y�����P�8Ea�D��D;�f��Kf�瓦�`+���8�Q�'�(��\�{�-��='�2�p��c+��Bm&�y\��h��!�kv�#(���d#�g�(Z�T"MP$!��D` �'�'Pk7�����;�5���voz�د�i�x
>�_.xۗ�n���k���p)L�d���h�d!C_) X�rMl?���|����GڷLȇZ �t�U�-h�C�c�J��?�v��T4!��;���t�h��׼�d��>A��Ҧi����Z��|�(b�^1N(�c P�l���x1H�h�%t7Q���L��|�7p�Y:QO��(��'o��N�l�詨������������)���b�HTGw�� ��2٨``0:�Ҁ9y��FM��U�䔓�.��|n��6�S�����aT�#WЯ��c��n�"� �z�4��4�������ѳ�G
U.vN���4uP {�=�Y����� �%�/z����i6�����;W�,k�������>f!c�OC�2�b�U<:^F�N��0L���kp�����7hm0��cw��=��և�厖!�M�����ơ��`�����}�� $��w0x�|��N�)nD�3�:��a���$����W
m �I�����f�P���ѩ����L�H���!� K�^I5�;㴃�Ί�����j�ˍ�P������������W����g>,X3'b��EQ��ƈT�=�T��[�4?m����Hg�6D$>�Zi\6�c����O�Ð���WM�-�T�T�֊��%u2�I�������/���h�k8��������+`V�ó{�i�����M����ȗ�^8&[��m��XFEFX��eݖ� ڈV �S`e0=5I3$OW/p��~�1�VԜFX%=.��k��Tı��s��}C�TS3�1��|V��x� �6�?� �y��-g����V��">4\Yn�w��řI�VoN�Ә��G���ޢ��\��֭�a���zGЍRc���%r��h+�J>���9��`$w�_f�*�T]�A��[n��bR)+��Y�G ������[&Aa0�XN�ɧ���OXB��$��BȾ>��0�fΝ+���j)܂;h�n�5�x?��Cu�ܨ�5V�0���jg �/��ohy�?�';]��e�S׺�`L���:�!c_�f�=�+���a��N4�~w,�-ڗ���S��C<�m���,_��X&'�g��ݠ��Q�m����B�J��L��t�h*lMTș|��S0�+|=&�Q�d�y�B�yY�Щ�6t�Py�=���U��UK��]e2�@�S*�nT�Y���:b@�B���ɏ���ҝ�� �ԟr��%أ�@�?�q��}1����c |��\�8��Mٴퟴ[���&w��h9e�<�C�k's�;�%V�s;��W�d�r�4-WB@[������J��g�,U��m�E!gNH�ߙq}C+��fyD���y�4j|~�����.Ɉ����NP����l���+T9'�Az|�nj2k�?�!e�$.%���*�e}����W�"<�Y�_P~e��Ɵ�/�(��m�1k�c�2��.�u�:|� �|~T�
on��4J���!p����ܵC�_�{�S�� �^��$,�����۾����RU����6�K�~&D������P�	.����L�R�Í�/'Z��CX�8���ҿ��l*�sI%@���锪=�X��J6X��������V"�����?ڤ�qe��������x�=\8���pf��0�/�~�>Z�~!���ը�B���"-��)�1*J��I��3YB��e���8M�ދ�R.Wޅ��b���kvD�#���j9�k>�?k��I��6��m�Z
'�r�\����O/��=���E22d�sȕ�ў�bs��<�S+�?Ec�d�W�vu1���/j�N�zv��y�!zcew�O?g�b�*���[�t��ٓ���S���5
4d[�85i�WϚ�,������GSL� ��K2q��g���>�sq�9|h���3�)���'$"A�p���T?s��C ي�/,ugn����I�7��e���e�U�mr^p��Z�n��8a��~�
�X%ӁJ���bG�^t��c f�o�j�f�����uX��ޜ9T��R(X�N��Bz�F��������l��Q�:�
^�	��&�����^NU� �L�4�V��@B1Fo.~9&� %�z��L��.<Η�������Ȕmd0�&���,S�(]^�����V����A��3[$oe�Jæ�%(|�@�}j%�;�c΂�
�� �i�ް��j����*�J]NsD�\ ӗ�o���4)Č�:SR�M�NZO�lO��jv���a��.��qI�����:��X�4Q��.K��zEO�y4��u�!.����Źѽ�p�?�H�	ƾ�%����9�.�.�AE�ʵ牄ޭ�{/a�T}�媐H\��Ė��=.H���+�4|���;��Ӄo1GR3m��)�l���CN͡��4�v�Ɖž�vg�\��t�>�d�����y�9N�����-Z�PU�qɈ��wI̴A�ʖ�ɲjX�nt�A���I}(��<�h�[�'j�Ӌ=ӣ���\V�]��cn�.3�qZ�G��bW--J�b�^*0_�L^b]��q,f�i�:��)��,VmN��ë�d�g��H�:��ڢ��@�cP��4u�J����A�)Z"����s���Fߓ�T++hS���;�nC�@Y�*Ow��4�����.7b��!Y���UfA2�Ą�=�.��͜xJR�I�h�1%�8�h��������#�ʿ�L�}Ȧ�G	�o-ME;0⩨��!W�q�at�r?�ΟE�J\D��6�R8J]�Ƨ.�AI�\p�ȓlY�Q1�Y���8�˝�I��g�<��o-p��W���e���b���6�_���G���_4�춰��Zy�G����c�����酒}EY1�Hhr8��I�S���%k��t� �0=��=����w�A��Ԯ)�A��X���N����\���G���e��"?Φ��SX���wF�N.��X����lS����B�oܽ{�n��L��SVɬ ���~�a����Y��]�x�7�����Ϯ���kdn��SAB�ܤ�q���*,�q
6�x���~�~���Փ��Ȑ�Q��!�Ns�!�t>��h&F�rǔ�ܷ�b>;��I�X����J�N$vf/a�gN=�fv���k�˫�wi�A�Z��s/��a������˷�߻�
������SW=��(�=ϩ߼"�9X�m���+fj�-!��%�""|i���*��Ky�H+7�.e��m��Қ�]IZ�$@D5�U�����
�sfm����5��_B�8zT�g=N�]VQ�-���pY`���p\MU!\����k����<�'� ��
�@�v��C�ƶ���j��VAu�t��Q��.7�\2����d�o Q�E�ps�����4w�;���?t�\I��%�oA:��$-d��@�A��@ƣk�K2RAU$ >�D�k��i����C۷��mW>nǚI�|���'g�3��5����N���1^��vz�ۭ'~�Pb.4�v�_VOGoS9�*C �9�1=���D��ˋ��[-��6�v� ��ɲ��jB��Z��F�����I�)��Q�cZ�9M��1�x蠛6��l��Ueco�l�Jq�ͩ�����NC��xv!�8�vEǒ�v/U����)���J���CO��\3q+eq)�(��UhHN\�:W�\3���N3���b�E�kPK�1cc��e�;����b�3%.�YU3A��U�� 
�~�w�*��9��.QU���T�1� �e�K�%^¼
�UmIJ��&��g{|��b��8=��d�_ u�t��[5�1�_��ʤ�̞k���9�����	���lu�?D�`��"Cѫص\̧po%�r=�����F�yc��V#?�G��5&A�*a�Q��
o!g�P!�ѭ1#���#cX���WI`e���Z��W�]/|D1�r"��&��)�&?D��T~�6�Dc�t�0�K�|1T�4wA�ӥ3yS�[N�O��N|݆~��F�&h�#[9��
u�(vLAm72��:p�fW���m��L�k9�������JL�:��6��G��]w�����!�[�&g,ĉ�+����"6��J,�YO�k�[e`��ґ�� K����Ċ:j���4�[�w���v��*�.@�Kg����Ο�J������=�Ǥϼ���8��K*F�)Q���P�����i��p�!ּ���숞��c���CY2P("�)��MV��� YԜ�'e�${�'�k���:��7��d<�5Ƞ�iwu��/��}<����R���Ѕ���A@S�!�������X ����Ľ�YZ`����U�IN�rE���O�/��׷��x/�7YY�o�������ɷ��d������6�GQE4?��q��;�BQ!��3xb=�����|�n!�ܻ���m)��)�	�|�肈2���Q�q}Z�$�:�M��<+��/l�/USNj¯�ʥ�y�~���b3.���v�Ec��J��]���2���'��q��J�2�����Q�2i�+b���~��}��X�4
.����8���j��-�,���QwN��\PkX�ꭤ#u[��`3�[��nY��j���/�h/��R9�&�{�\[2qX�UL��&�$v��H�Q�U�с�8A�q��vN��sP����&2s��dg|�"�T�n��kl��%!lGc��G�e���ۚi ]8?�Ux(4�ab+��'���8�z@��G�^z+*����\:l��)���)G����+�*2IW.��
�u��t�o�It�s��&��N���<��?m���� �'8w��|���>��(&?b˜����S�Jud'��1z�ݤ%�'|Ly�,c�'F��Y4�%�Eg�*6�{��s:vyt6:!���jqDd/����u�X�ʹq��,4�-�s��6h!~�da�s�G?Gs��-�U<�b����~l�u���6�R��0���L�5Rՙ�l�"� Z�� �;�B�|j��4�c1�O�Y�=š!�aj����#|��#8lH���E�|��������3+�}'�E��W��	p�pg�P>�M:�"�YIp&�����#��&�'E=��!$���}'���������|U5��Y���Z����Y��kdG�`��Z�wؾG0����_�fu�Q�R<�h�������0����M�}9�U�(��.H��5�*Tf��D��Z9gRmF��w�t,U� �`��ݮ���-4��'������8�l��iS�ɒ��V�G��	�+�*�&{�N�kӄ؜����whnH��ҝ�HS5�~n����3:�`}�@����{2T������|F��lpUz7����.eL���t;FT�^���\MH�ik"t:,���?�3��b(~�ַ�|#t�����[�.y6_�Z9�~��	T�3z�N��R��~ k��Z� 4>�h��q����`�\�0�����y�_7�~ȫ>_�QM=>,ڿ��_VMY��}V��ǋ^+�Ihu��E~$�]�3�d|}��W=�`1�hzu���"'恥
y`�f�CeH1FO��У��o$2U���t+ʏ�;��lǄ5�u�u�Q֣.�A2�?6WD�M�������܈&��������V�����#P�})�I��@zl���~�^C�o�rʴ�)H��,Bxe����r�U���[w��l!=�J��3E��ҏ���23��|U�8���(����������1ᓦE������YBn��-�=�([ժ��kwM��|R"=�KDnV�Cަ�6����閾�Fu���1\�َ��=_��LT�_]n���)$�V]��IpM�i�ě'׻(M�Ļ-x�����_��E���;t%��5��
w�cB��1�ő��Y�g�L����*�I�h޴$�S��q֥������UQw��!��$yz�����((�<���a�q�L|�a���q��S
ϞE�B�%�h�?J]&�(�X�S\���&�j����c��֜o`Bp,]Ě�v9�	���Y݄�+սj*���sh��Q�ź�vC�����'��D9�L�&{���T5�d�F�ڼ�'r_I���A�!ב�U�L�,L�l�l�(��*xr8(�ck���?º���PZ�.�&�㴅�ٲ?Ū�9W��1��_�]���VP�Ă��4���k�Ψ!j���X6���` ��Xvz��	�~;";C�C�0z��V�+�a�֨(,(����|�F�jbG�`M����H�����I��疲���@E#�A�
���X�	S��!�cWO�28�����j�(��r�^��E��ō6���{Xz���`��h�-������d��@'c^�dp ��ۗ#�l�R����"K=��Ns�*��!T�܏�I���SY�ܥkw�&�+8�'�Ԏ�"�����+�ȣh�C���r�4�%y�]�J	I+o�
��2�%Es��6lTf;`�EO)i��������X��iH���B묯k�.�k�7%��p�t��O@�� �3t�<�u�ی�b5?�u�#�K�!���P���Lx�[I�b�(�p�S���di�B����y,K��:X����/�<;\N���j^�Z.ӿ �F����u/�dT#Z9�2gV��l�d2�/���C5P����+ٲo�m�ǚmR��'4�~��+h.��1($!����=�ⅨG\Q�~�<�=�����dlp_�V��DJ��O���|����z�F7�0aU}c�L`A�V#�Xi���$$�Ţa�BU(�M{��-��A/".	���� ���=�}j���e Cv��5����$똻Q�m�=uP>�6<�ݜ؂V�������V���.���v2~ç�̆���O9��K;�DRw����2''���ݝmM��J&r�[�?�&$z*��ՠ�n����ĕ%�]�{)<�$����������� �����z�**o�5}_����e��7-�@33��J���/��5�M�t�%��PO˹��mM��c�`�6�g~R)�bG]q�t��
�ji=߳�^�)�²�x�]��kZ��a<�^�^�7/���)Q\R�^��62��V����Ɓ�` �z��M^!�@��~��Hr;�u��C9k�6�xY�5h� �^����F���D� ����q�dJ;���ϥn�G�5[�A���ñ��'�К�MLDE��N��H%�RƩ��GEV�Y5}��;�������H��a�}�qM�|pa�}YJ����J�-u�KL�V"F(��w߫��*�JE�����@+�o��L��l)��I�(Xd:�N���Cuڬ;�g�3�U�)��b>���^b�K�(��H�K�I�G6��O�T_BFp�)Gt�]:�:;X��cg�U$�.��|e�bĐ���$�x{ �W�B��P&}Ɣ�(��_g�ë	(���r�����Fκ�1w-;˫+��%�鉢�n����{�N#�oo~�r�S��U�o�;��{��#���V���&�G���>4���t!8��P����D��-�XP��v��~�%9����b�&7(��?(�8��j@����ꋡp��[бZ�M#�!ʤ�1Ǥ]��7}�ӹ� k3TN]h}%��w4����蒭ճ.�Jv�;��O�jN�'���;���mJ�	�������l'��]~�F�گ�]a�]{2wY�"��`�&��C@M��z��������;%)H"+Qk+J��)L$�TL\����Y�H���0�vȷ��7|^k��u(!\����r6mbXt�6+v�hZ�ڳ�!�iž��v���jY�L�S�kby/p��ʵ���u�I[�	�%qH &�a�[u��͌���-S�1I��P��ue.Q&踊y����:òSi�ڬ�2=
|֑J#ַd�,�B*H�"vƾ������f���`���3i��(H��QVq���}xZ�%t�K�N��yx��U�8��r9�_~�=t�͆�F��'�Q-<0���E�G >/�[ ���]^Ԯ�C��&����)�hs�@O�o�������ӲO
3� |�yO�T2�FS����ZW��S5���3|}9�eH��.y#)���{����:�;�k�2����-�/�'G����@M�Y+� [ ����	�2,JiԍF�俆V�|̓.��9�{��Ū1l���w��܍Y�����Sv�/��WIq`x��:��Ҵ� ��"��J�<b~t��Ռ@xL���Gn�'������8�����*n���W�E���B@&�՘6]F��̃�OsѮ�C֞w.��L>�6	��ܗ�'֗��������Z.�f�af�5<�5�>6 䢩 J���:�؉��.\�[���_����X��tӕ��zU�Bs)��1n���ߩ�+n��b^'x9�ڌ���W�XhꆋPe0���wѼ�}���.����F���B 9�����jq~cE��V����S�D��{���@�솒Z�=�1/ɵh &�)�͠ế��!�26��5�ꁆ!n���`�d\)�}pm���m�qW�k� ��5�+}�������Y�_����>y�d^N�e�44�rI��:,I;t@���Rxs'A`hd�IS#
�~�ԛ@�N��̄Z ʜ�>YzV�3�7<�q��3?*��#�w��d�h�nWL��XX(�8�U�$���Κ{�����ҏq�q5���Tn�\`W}i9��/\2���q0��$؟�_X�* ��B��} R+���]కв��7q�*/SzMЅKkEB���i�&>���`������Ӹi�G��Ɔ>Ê�C�=��iI5�1s�6?,Я�y;�����&@!� ������XP_~���Gz���x��S��ѡx���v7nN9���jQ��;abώ����s�W䦵ɵŽ��L��S>v��v@oY��6�ݭ���$��ʍ���n�Ϗ&�࣐�@�Y���r�sǺK9"|��dMeK�S6���_��LO�(�n�k��%�D����1&�#,_R�^'۞�8���Id"�����|}�+)�4����*y�O�hp͉��f�T�j�:�����H��N��g�ϥ���v��u��!�æ?��vbjf�+�Ґ��o�.����������i�<�4�ƺ�/A� �1��|�+UWB8 �� }}]�7E�C-F�g�`��^���Cn�|>st���zs����|rj���u�1D��8�ُ���/����V��-���\�9���C޸�dۊ�_�¶�J����a(�q����m[/�R%����Eg�����͐�شT8��$��SǨu�h���g��M��T��5��u���g�6VI��?�N�[۳P��"�6��[|�m7��88c]cv��Y���s$����!�}uM���	�ɿ�QL����<<��#ʪ����\�w�-� ݲ�]��)C?������]6vG�ZƘ�-J(Q��;�	9{��k?���[��'p,�H�I�7ME�/7܁&��I�	X�@��2(d*L��Ŏ��'8Fh�¨Ij�-=�M��=�y�mQ�&R"��M��ai"nP�,[�nI!�\��]��<6ԯ���@�ػ���(��:���]�h&ԏ��34�q#p�Tu�{���v���^X�SG�3YEaQ8 1�~D��v�ޝ7c���:�	���<�bj���t=�p4RT�/��c�Dw��kAЌ�P�$���*4�}����3ȗ��vhW���4Mf����I%ų�\x�PiD�D%_�}�Q��йi?��W�A���Bg���x,�g�3�:�t1����)S;������!0��ǋ���h�v���X�X���+e{~j�%������$�m��=�jD�����?��4��(�%`C��M�cQ��V�zUчU���D~$r�����̾!�;eH��4$}�Q^Z6G�e�o����c�HKf��Z��uP>��ݭW}4Z��O stc��0�U	���T�Zݕf�҈G$�+�{�-��I�/�0�n<��תR���A����g�K���O{ 03V���4�ѕ��kE�]�_�����f�?�䫨٦��R�����H@QX_)�H���R��&��v"�4��}�H.j�����l�zye�Z���IOk'
sc\�[��w�wx����pצ�;{n>�<�c)ҍ4?�P��8|{���g]��r��F�!�Pu��&�����1�|>`�YS�^ǈ}��H5/�_�IS�BRh��G�;���6��敾��t��I[�AYw� ��-��&�U6�ٜP��v����h��@��!����7"�����ny�K���D�{.��o��?�.Eŷ;��|J��d�ū�'>Y��	�����I"��^QGQܬ�"j���?�C�X�q�M V�`�&��(9��7��-yXMt�I�L����o��%��/z���lh@�^�:?���)���`>�KEO������D%s1f;����	d$��L�n<�<*�$�u�,�7�cj$���e�*B�#݈�|�W$�Xäy^38i�{$[o��T�G7���lTA�I_�����+��6 +j���;�Q��V��]d���g�!�2X�6K�72����Mh�q"���+f���_4�<�ޥ쿀]'|�vP6K�\5_�Ϫ}�B�'���
ܩ�I(��f�y��ܾ�A�LB�rMR_��2+�?R�7�&Z���u�GN�kM��WK}�[t����w����>շ�?�ԧ8K���hh�򖭮]��y�����K������o}��c�5��uk*5qQ�ԅ��e|1���xO�q,����<�C�@�'u��|�8����x����;�[�2�D�PV���h�"�mub���m'*� io����p��w���?J��W�Tf��#�&-'�s�����3��:�ٌy��8>�
��Qv:ca�'cLƥ]�]r�yrG6�d-���m���P7gd`Fx� �"��n6&�4N���L��Q���]<<��T/��c?c�;���$?�^kMFA��I�T� g���M���Zg�� �	bZM�	��LHC���I��38�?���X�DԶ%��������u�e�*S.���+8ŵ���h �˴Q�)�*?#�GÍ��-7Bt
�X�W眣����Mm+.���SN W`¢3G������:V�H �{	E��T5���L	y���r��
s�j�i��I�Ac����-�!��H,^�<�'���I��y��l5�k¤��,��,��ߢ�A�O;�@
��d�Q%_H�P�y����v
)�K��j�!�����$��$������ �+��E�D߉cw/�t�����a>��7x�D��@��u��zU��&a������)����=�P|_�$��o%�|���d_���u�x��\� �/(/9��=8 �CM�Z&���T(��]#ٯ��r�+Ţx�56yov
N0]�z��j��w�h������i;F�TC����ӱ���)�F����"[�&'��{����Z�����{׍۩��Ւ��7�Ww���b$���Ju,0���O9Os�N��;Dˎt����*�̊�R��)[�Q��k柌�z����
�bٷ��zFkX����^�D�d�v*�1TV�#{<\&C����A��'&�9+�~�j7F�1ɡ#{�:�H�v��*���.�c��h���oP�;�JF
^���H:z:N�E���oZ�s���qKҠg50U|o�*�v���~�ڛ��m�+!OK�;�#�4��L�"�7�
�DbJ|'�T_�E^�m��:2�]���i�̷�R1#��I�����L�^��-�F�NIiԋ��+#h�R�	c��_�X��J��Y,z�#��Q�k'cȃ���G�s#��}cY��#�uڼ��@���͵��&�~b��쀭9+��R�'��)�E��m铿����J!���Z����2�I����a���
�t�k_bX���v���Sug��@ڟᵵ(��m���v����hFNS�?mu#>(��r���(��<f�P�p�k�C�*R��D\e��E:%�נy�Bf�p<B��5�A\ l#)�v�N�77އ��lA'ES8U7���.��?��a�0�H����c$�	��JBy2�b��u�p�yh�rd��RN����ugn�v�kh���bH���b��ɦ�5]	�bC�U�����s���c���0�)Ï��c�����b/Ѱ(\�� 툢�F�8��^��]��s{RK���?�l�r=��s`;�&$����M�$�6��q�Q;׿3n�Wr� �'0�d��+�����i6�+�+�dV�mB�O+b=GV��=,x�J�-�j���bi=%RY�;�>�����)�z�䬨����:�%G�m��C�x�j
t���Qf`�A!*��g��f�D�Ӏ�"�ֻ2��v��0���o�8f�Jf(��N'�Os´f�c|`��t���bd�6�[���c��A�A��:U�'���s��2���� ���ϯ=Q���$3w(6I����q�1l�s	�n�yH�.���Eu��(V�e��nK�`a#�R���[2vV�t������DLp�~��)�����٭&`2*��o�@`v*�&�G�<)#B��#`{�"�q9�$a_���W �H�
�E6�ׯ� �vx�s�u�Ȱ��"�"�[�؃�E�1����XO*��\2�ud(�+"v��#�d�fٰc��a��WZ�2���+]@D`��k��qqK�ez�����!E�o�}9n
|P���X��
�O���.��n��
��Դ�Z��(�g�������'�{i�4oi���~.B��7�#�V_)g�-�#���I�>iB��{���*m&Щ<���A~�%��S�A����[!����Aks��_�m���ߕD��N�8`�z�0�p�������^��D��ʢY�|�k�-̉���jOZ둟.W��"�4�]�����d �����v��R;R"&1)�3��h)��(���(���؂��W$����U{	��%�7[������T����Lj%{$ٽ8\m�W�J��u}Re�0lv��� ��J��&�]��D�UD�8n�6/������Xl���l6}`ʨ�^=�WʃA����w�)h�a��˓,���Y�p��C0ۥ�Oa&�r*����4������5��g��8 �W���f�wO\�ym4UW�ޙyhS����~8N�j	��
pA�3m�~��g^������h������m�4T����Q�����(e��0/E(y�j6�_)���!5b�eN`uW��eƇC���a7ޚ6�#&��_MHȓ
�x�
�B�za��5�φ��C�����<��#D;����!c."���7��� �j���yGÚ�B}�=�_��tnНhEY:�5=��q*�6"l%L���8b���zyI���J�x:���o�,�5�h����#�p��DE�Ն�~2E��4�v�i��l���t��9xC ^T�|"vT��9Q3ԙ��F��$
:c4�a��d�/��I��薒���V�Š�P�g��t1�"�5����-�ޘ�֢-wb��d��$�f�p�~�#��En�.v'�O�ޜ��D��&�`��dn)�BxM��J� XŸ�c@�KC��g�]w��X�|�ڙ
��m��C=�,&3��H�[�w��;��Κ����Imv%\/���o��K3�haK�K��{�|L�ƯЧ`0���|Zk�H�x����it�3��e�����3Ր�!v���\�T��B����6�!o��dHv����n6���c���F��Cf�I�,����YԴ�.�W5
 a5j/��S>���ɿP��E,��._��[�FPC�jm�l���iW���J��3s�#��d^���mв�J�<i��jU��	*�DkA=�N�0�=X�~��>=]�����9�'`�3��&P�?��w<'�����&�]ӫ͵�J��b���L֋޼�*�l"�dT��[c�C���:5z��Q�B�k�꼟0D���tk9��K�U�lŧ4ao�|���v����z��˗:]���M)��B���,����>|$��&�g�ۥ��,h��0L:L���\�m���B�������9/�=�w���f��x�7b��{^�)m��\�]�b��>�s�[փ��#��0�#��D
��O"Λ�'�(�x(>c���D�Qn�g�si�퓑9���� �{����Z�(BzR�j}��VK$d;�6�텠�l���T��5�~a�Rđ� *_0%���\K��Wa���:����D4�﹑���N.��md� \�A�i-�MR*�W��f����G����~IX?L96�Ɵp;+]1��rm��.{g����W��bě���ph���~�[r�Q��:#z�{Ib��[�|����3X�Ig��un�;Ft!7w�����MʨǗgS��{]����CV�X��P��">��oA���K�;�Ҝ��}R�sJ����m��f2{S�V�7��&ؼ4�j\��;����x�&�M�i�e���q�e��gmp(G;H��;z�������By�=4=a��[�j��}��J�|ܽQ1�����Ap��νe���ԃ*�bo���\�.E0���>��F:'��Ҏ|��?
_9L��=��hnE`���h�|���T;)�Cg/4=��r?@p;��� ��2Ӄ�����g~�ZOR���� �H,�lL�@�qo��fܬ����}���A,X�$�юb4�*��~���0z!Ӭ#���2��VR\��u^?#2b�p)��z1~�����I*8Y�k�o���T�i[t�#sbȞ��|�����P�7�.���6X�����,-�ǀ�	�/`���l�ק��/������Fͼ
�H)OA�z��?�!���轙­�%t/R=c*��r9�cj��3U��ٌ<�$��ɫǽ�J��nh9����W�NE�� F$뷿㦻��<�(����cPO�s��󑏁k�j�9@d��pg�MhR������p.g�=1�P��{�*!����-O��݃}�&����YW���ςg�j.��@�D
t�qx����J��N�q����}A�D�3��b�g�I/�?�E�Iӆ�>zX�i8),�5]�VeWbVǪu�^��O3쇶!��x��|�L4�_AάW �:�C�hW�ߌ�)���K��X�$���,��Ɇ�f�Ź\�vL����
���x��A�u��2`��ӌ���������>����I Ƥ���װ'����k&�x�2�_�l�ꀐeQ��.��5�񌕋`ywJ���e1�RR�/{Z��� (8
�F���!�l��5�F��0�����pl.�x�lʌD�N#hHh{HG�A=�:�� 	�������L�:+��>f����9d5����T��"�c��}����i������64��,�Ug��z㊆�J)4��=A�ƴC���V�U��R5���u��^UV�ԣ�2kK��4 v�w�j@G(�����TMЁp�0T�oh������nփ$��PX���m�A��ki��[��,��m1���ȾM`;�@r_��ԊH#����UP�^���e`T��m��ǧ�n�A�̦��nB�����L_�����,�B�S����FOC'���N�87w/��S/�:nr��[�X~�k�����ţ:͠��r��r�tD�>�]o�J�����G�LȻ���b�����i ��S��㠩��@���y�AD���X0��L�g��.o{�*cإ��(Q��Sr��[�X����5��)5���#+���
ɞ�⣒�)�d�������BT��~�}��^�?��Y��)�t�e2Okܪ���
��g�x��h�^ ��ف��v�ָ�-5�t�M��ͨ��R���nA�_��Zn��L�t�l"$�>���C�!�q��_b�/9f(����gf�#E ��e%_#�<��"^'�K�^>n3��]�+p�?���C�E(F�݋�S�/:IJ�%�<dTsi2��_�j8�������s,S
�5��F���ʛ���x�X%%kH��ˠu:���x��6�o{����T)�Q�v���Ѧ��ŸZ6�zp��< |��'����C�ߙe\�y�T;����Ho�J!U�g(�u��cf�o3���E�:a&��|�����3n}}����X�R�~:Q=����f��qu���37!C6'=���p��T[Ì�d!.��P���2�{���-ئ�IX�6���@�{G��z�yYef�_LOq|0��@��f#�pV]�:����be�d]����L�H����)�Z^ct��'vY�)�0�Bk�]g�;�~7��V�u��X���J�(\��,�_E &�4�+�lA=/�#W��l�F��y�K���ҭ���P��!y?!�t���]h�X�{�A#w��7�G�s.�Y�阊��� � )�9Q|Ӏ�L�(��>��XV���p5Bk�$�`�;=�j��}��H��G�����m���J������w�Q֊bv�/�f�2s/����h��f��4�6;}�o~=����<P��N���]�DM��a�i��!\Gf��J?1�r�<áL��f�0���䲊N!(n��?!��yx�*.>=q:r��������4��j�e��z=�����D_����^'M����<��TLx�H<�nGժ�5�� �J	(αA�#�����2k���0�u>?����9�����N��q�s�c���oy&�M���Kl��srL��t�@$�4�W�Qx��3�f(3f�l� �G]Uߦ(���:��Z�fcq�U{����o�L������;Y��V�
��)�v�-.F8�M$�W�l�>��G�$X���@�<�<gx�M���ϭ�H�*��Ty睦$�����Jh�)�l��k����jI/F�T��G˟�	p6�2���:�D�?x�_&�J��/�\=���t]A!����~M��a�7�܃�.�E�������+͌���"7ֳ����ĻS��%�n��d3�~�:���Z��\>i1���ڥ���}j�Y1Ƶ�q�H�������p�_=��3~���PI�c�C���(c��I���5F���"�#l��&��b9�k��*1��#�ڷ���s�jGIy�y�S���	�q  R�f�L�Ρ��u�e"/�v2�O���i�Q�3/��G�}-��u!?�ΜTk,��~��W�`����b�b � lx�,`|�����?74�/Ϟyw	�Ўƥ�����@���3!ʕ��Ҭ��H��A�,��ԙlA,��̘B�K�#���H���*�х�H�K&Sȁ��mO�c�6h{������KO�s�.�5��H-�۟㛾�������3����"��"<GJa�g�1�Yn�%X8�@�H���j�?f�B��E��
`�#������FQ[���k͜���3�YyJ�ɚ�,�Y����ea�g�A1�F�A/�.i�
?��ԮpJt)a(Cw�k b�����'$�X�u��2�gq�D+Z]������e/��$��8�2�M��|�s(��a1�3�Gn����,�J���%.�x5:<�Y�ev��G�R⋥��k7~�>�C���Hf������q�}H�M��
8}��|Ga ���7Q�}%P�$.�d)�혏�o4Zh|�
=�xN9�
aii��(�<u */`Zp��������7JK��9�+ڣ��-�$6��t�ѥ�$e��B��b�6��)��BS�N`���8-O���R�@Ѝ��v�j�`��������E���c���Z����]�@E�I�w�������U�s&I#B]u#@����U[���8A��B���&I�݀���B�b�|����sp<��M6��C0]�������eC��c�vsZ�Y'
�k�J��ؘ~?}&��u�<mGA<�;����pG�pp$㜮&�'��w����tw�˂���1Bbɇ��Ϙ�(4������攦PrI�p'h[���¯Z���}�bQ��ߢ�-�mK�l�$΢f7�pg(��S3�{޼i��Rv�p2��
�S�}ֱގC�Q�R�N��[ש�|�"��|�՝?�xɎ�y�g(VE��T���R��On��&��M�P�����Ʊ++�<��<M�fk�Q�>W��R�#��9�W��c4�&pn����㛐�]m�@[v�۳g�`����ބN����f��m4�p��Q���TUM�M@��S~�db%�.�%b1"kQ'O�֘��*�+���P�� 6�
9,<����uQ&���i�*���C�(<r����[e�Ċ���)�-p���䏌~Q������Q��Ϙjg./W�	�UY�}�&�T��~�#���q��ֶ�	�}�J���ni���/Dy���{J�FOx��u��F�F>���"f[�ǰ�ns[^��͊C��z�5��wDHu�y��t�F;�U���we��_͟�� ���-F�&�jD�ub�Q?�R�k�Կ���<��.���9荠�ok�Ed�z$߇dm��́C'pа��-�O��� �&D�B�ʱ�Uu��9r����>��d��� �.)�۵��g()����=��l���^|"���K헯�7']g�[WZ�����������~�J���mb`��2f��$�P�*�C}�ߦ�����Z��{����R�
�k0w4�Ā�S�MQ8Cf�;nB� �;	r�MX�a7��Kr1옱�X
@{(1çb~�;>m5�u���)L�@�s�7_J����`�:���+�0H�;�{
P���m}Q��`�w�İ�Nu{�j��i�p. �)�֋B9^��Z���U>ģA�>%7��Γȼ���E"Ej�!�#���+�oz�ej���ՏH0!�f)9�̅R���E���ɞ�:ł��1Dr�i�[�:�N?�l~i�ЧY+dWV�w��GM�f�wŻ�Ȩ�S��	+ޭ�|܍��
O]�k}��t*@�TB�u����og�Q3g'֋���G�d�9Y�����������}�7�^b��Ɵ|}����x���J�-0.R��v�-@sL �!��%��, �
��Y�ShưJ�k��&P�Jm᷵�d�b�S����]0��wCbW�s9��}�@b�6a:\��m�9����"�P�e,���qqI]��_�Tl���_G���Y��HT�F�h],"J~���M�~J�SDULS�n�V�q�5C���^2��z��!�`C�/Rǽ6���W�x�cE�(�����u���f���'r�0�o�V{���+�Ce��s�,�8\��cr�oM��~ޙ,��ӕ���y��ng� sQ�/N�E�Aq�P�������cpc�[U��yr�ʵ��\ǕD	�kkO��E��<N��e�@ �ӂ�I@-ns�&�cvP��Z1n0]���	�'|�[	�m��eF5� u��t���T���(���Þ_a��̰Y߫q���}#讝��މn���dz鴔��6�^"{�aKm�}�<2�o���u5\Y�F��;��(�b�c�6�i�;�]������K��nt}\��w�&���:u<؈p�.lģ��������)�������cP�?I8"lD�y��	�ѵ�/g���4;��2�у�{���'�/��Sٯ���W�`8A�K��0����K�6]$�����x]�������6[���ڏ!&���5)]�@�q*-3����tʸw��qt��[3��\���H�W^�X�7em�x��z��p��;�9��w^�Z+ݹ���˘�d����Q���]V_"��S�q�rL�.ޜ�|^>{�,}��e��2p�z8e�2=��U|9��� �FU�u*uJI&x<̎أ��������:�A"|g�Q֞dqG��w=M?\�.Q%��j�����3D4#�qds�ak��-��)��`mȎZ<Ϯ=�]��$n�
(�o
(R͸<�~:�a���u1@A΄��t:�z� �hWE�`�C;6��9F�ͫ���D�9��G�t\-R{?1kW���r�!��}�#��àx��G��s��whs��2iE�8���e���щ7�*%%�ri(�Uno^�B����م�NH�;n�G�b���Ev~o�g5h(��<�� �Ȯ{Wh��
���?.�C���^ɬ���!ߖ}�^d<���ع��~����BG�{�1t�ׯ�����X���U�"��2�O���Y]ƪ+����$�1�׬���-LK�w�K��-�{2��P�Eny������6)��B�*�
^�n��k�����B�F���e�8������/� o����1^���Y?�6�b�n��˞}�u������{d� R׉D8�'|`M[�0�������6��N�R���9?~z���YS��l��Ƒ����by�<5$G���ܓ��l�HFU����а(ip�#����b=�_}�� �PC�hf�5����g.��e�u�m�#wQ�:��r�Իׇ�?��0d��t
�ᔪc`�v="EA���� <������5цi�[Yr�xbE��A�¯šX��S$������r�#E�r.�T��im�>:��>�������y�����2�@�k�Z�o-��Ց��a�� 9��2ǒ&��6=����gH��p�tZ�^|�D������'E�s5f�+Vǈ��;���cQ@��e
�PP��9L�z�و�n������h@�
Bս�O�<��������@��V�;1�x�
¡ gd�s��1����ER*�g�K2ېUyh�j�:�q��c��lu�X3$�v�B�)�*y�����M=�v�j��7��s�v�eho�}�����������3/k�Fb�1��/Nġ�X��v����D���V�7�k���褬����C2��a�����.�H/�c:	D%ֲG(�q[��:��(T�X�@�Þ��8�ݬ	*K�K]�z�8�"�T�3�m�/ݦ�;�����&T�+K;%5�%��R��$.%��"!M�g\�l(�VǞ�M��:�&�G�n h�d�ӹ"T�������KH���d�F�b�o�/���Z?9����G��V����v�n�!�ڰu�͖ޟ�})�7'��;�aZ�|��0T���्d�S��hNj�^���J���Vo�<ۼ��!!�'<8�� ��7wmj��hVh|�8[�?�E���,I7��ҥc8A�N5^��G�}%��O��}\-�G�9��ٝ�I���+��ް�~l+�iDG('�J���o���>��~��V-Ow�D6Q�U�Q͞�:���q�����m��;����XxV=6�J�/��?utKÀ���ɒzNIKkT(U��8���M8$4��^?B{5$��L��-�*��>���0k`S0�� ��|w��tn:ߺ��(	���	�E5~K���s�f��	�Fo�#=���H�h�̡&a�.����WuƖ���:���r���T4؃;)U[�i��v,�6ѡI��t0��ɀU=�k�=��v�q'+WohNn<�Ƽ���p}}7��Q�zQ� 8;��:�%ht#r�i��Q�))�t��~g�J5+i��8[%~U������VX��P=-&g�U�&l9{=^>t������Z��@X�Z^�Dk��I�פ��C�m0�)c�O���U7�V
9@L�O+���K��v��vDt��l�������Gg�hR�[���&��+�
Z��;����k�f	����>��r���),Ȃd�{|�.�F�9��C��2�U���G��?����_jL۴�j���� }4�c6j�N|�k��`J�3v�#Z��/Ka΃��M�! �֤E��������4����+��i���]K���7�r����7T�f���� (`OT�7x����xҖB���
�z���Ե&h8M˭Y�\�����<h@�:a�d�N�T��!E�0ҫ�6���7NQ:^�l�[D/�Ea{k��m�����x�h]��1�G9�>��� �S|G>x����۵��Ի��vA��1�O���{�δ���_E>����c��U�2me�&D�A�� 6�gN��?�,�^;���9��d�4�i������jLjq�)9��S*�jD� ��C�\ ?g'�i�ā04)���4�4�pB�R��� �r��w�w�a�.�=�![&��ß���+k���z�]�����x���_X�qb�?���9S�����+�Ep�<�ā��m��b>O�rCid̤ �>}9-�E���AY��<n؛Yda�a����{n��͆L1Gl�-ѹ��QJ5��!�F�K��A�\W�t��N���Q��3/o��v�T���h���鍓����̛���nl�<h�s��n�<��,���s 0}	s��A��{k\��o)�*Q��mBqJ���-���=d}ġ���A2Xyo�e�(V�*�6�BE����f:{L3Cl5-��b+?x�=���\r$��l[:����Y�t �چ�x���@��Y�G���\.�T>�d��m��3�V2�FU�g؅�+���V���(�pE�7����g�{d#��[b��2���LnΗ��.���u��/0���i�kh5�	r9�������}�Ud���ɬ+Y���B��/Z��nHF�˴^�\I��L߄�S�|t{��uv̌~ >�5wm9uZ���?����:
|�Q(����H/:�:J�C�6A�6�d� �-�j��^�<�| ��s���=���S���O���O���l/��xk�-^$�����1�j���s�?��U�\PA���U񹒌#����j�rh�-�dCq�8��?P����u0�wLH*�?��E���Sd$#���q)�;4��I ܕ~W?,[}tƄ�%�_��%�����߃}nO)�2WNM���x�]է#w[k�Q����b'��DX��ϟ.aoijX���#�=-�6��"h�+[��F�*ú�L�Z��x ^�"��u�<d�F��B��e�[$�d�&Cuf�����3QP�ԕr�K)��B!��IbH� �����L�0醣���_[�2���KE��ETp�7.]���ɀ��2j��N������PлXC�ٯ�T�GĲ��[��lͽ����>�ֽ����8��-n��7n�9O�m1�tu�n N5��4���L�	�Ps�:?�+L{�Z����� ?�-oo1PO��w�o�x��@J��ȡ�_vm\Dہ��\�5Q���$�=���n�����DPU�'.��TO{��WI��-
P�ݰ��G���GII̋���]V�J(ܾ�� �M��n#�:)(�;�;`��|����0����7�ͤ^�[����XOb
��3�?rL�l=�'|YLڮ4 �&�ܬ��R�Π�p�\�{�N�(l��"���SbIE:f��W��;�#�N��"���t�%2A������e��
�##%�|�ܸ
|�rB*�L�t䧏j �[���z�dB��5/??q�5�Z���G�x��e�>���9����Ya^V§��WL��ϻ�Ԍ�|�:�8�4i��KI��z4��4Q�^Y�������{7��Ǣ�ay&�4Q?��mI
�Et�X
:"g{��h��E��3�^ƺ�ժ�Ө�`�qr<0����dÈ�y�3nM���0}��-�ʲr,>�[�O�������Ű��W��.6��,j7�`��+�g�z�S�^�����Q+2p��V�m"^�3�\���ww���D*/�S�x�#���t�/� q'��4A�r ��Z���Bt?nrt&��s��p`L�2���F���-��9?�%�aǥk��c�V��}Jh�+5B��;~�{I�o�p\O9֖P`J��JJ�,N|��apF����)���'��M���rn�����i�T�QN�2��q�����D }�d��7����ypH���Ev8��iv�p�̗�K|]�a��Y�����[�87��7�E��70K05�;�;͍i�2y,��?5�,�tp
���t0��y��u�N	~��/a7c�`�)T�	���_�$�	��MҌ������:#�:;gv��6�L������*GN�ͤk[�UY�lŇ���pE�DvF�Z���x��Ő�W�-�3$t�U�Fӂ z*�����4���̔�x:��ix�V����)v�$���'��I�}���U�����=#oP�h{q��^U��$������R ��0���ĕ�	�?3<��v��7h�K��U*r�]�^����N԰Eq��6;V�kƗ�D�Y����6p�q���B���,���3���ê�e��!d�7= ��?��c4
x~���폎��R31�c8��"�#�j�.�]cb����[vf8[�|�;��ڜ�4#�ͫ>�2���֋άҸ	N�HS��q���sH�)��R����\a�"]ࡨS{�E��ܧ����>�Ɂ����R�%-�O),ņ]��L"�\4ب���Ǿ�x��'�5�����C3y�N�R��5v<(�HsX�P��jMV�����Ds� �Dm܎�mpt���l�"ʩ����*I��}���c��!�$e*DK��@A��XFf�FJ|l��-E�w���*�m�B�::[H�~�C�NV9��ҁ�U���ʧy��k��m6��(Z��P�}��lRJ=d���f��s~X�=�w�8ՉU�΅�y��'Ԩ � �����'q{��Cb_;��Y�B�-`TTm�	��1�X����w���<|j�~g;��b>p�M㻎%������+'#)�����������O֜��4,Oyw0�"��F�B�%r�2t�D���?I�HH�/�e��Nx"�`w䵍? ܿ��v����66CQz����y�G�nP\J�M��i�Q-y\*kq��E?LɁ�������3��l�I�Y�FT�/./�J��m�5kE�І�ҭ�}�扴?7��j���BL�4��(}x�w��<u��^����,4~�gv�+y����g"\��Oz7���i�5S�]%K��S�..�T��J�:���O�|y��"�D�4��9����8�h��8L��V�%�D�ұ1F�t��0�q��֕@���q�8�vbn�Վ�6F�t
��vP�B�~d;ǣ�Ķ�y5�r;���L*��&�g�*�3����v��t.�|��T��*���Ф�[2��`v�Yǡ���x�ԛW9���o`n�p�T�ￍ�fn���O�����5_�����V����5�#�!W(�`���
�̀ԟ5��hĿw����
�tu-M��x��6Ňq�,L�J�q}�/?���`��l7��3�/gcCʴ����2ّwsl�|lG���R$c��}�a�E��u�P�-Ȍ�_�h��
�{��%��V�uY�/���u;�q�U���.78"{��	���"��!�[sZ�IT��|0�ʀT�ƀD�B��].��m!5z��f�������ΐ#ڶ��GQ�[��f�C���L(�2$�܇��;-	V���IGX�/�[K/ݽ�ȹ� �R�]�!�H���1��
�Y�7�/i��n<�gf�H�ل�IyT�%��D\ЗA9�F������d��pMy km|�4�UN��pYά��A���3c�f�������ZcnP���m����D�=�ǰTOM,��S'%E��U�oGS_�{QW��J�U^y�?��A��86�(ѧ�wм�%�)��y�ԄZa�� ��Z��d9!g����0�u��q��� ��wg� �%�R�i^������Kw���ђ�w�.���*�����y�(_�G�ŷ����~Ը�u7�Yv&�ə.�ɬ����͛�t´�&�ِ�֐�������?-S�è���˪�;s�����PJ�E�	O��{e�";Hw\�,��a�q�m� �$D�$��"RgV=�0��r�Z)�2�� 8��	.B3�~�8�.����g�0.�{�f�4��'>�R��i
����qd��w�1���\�=����'_�r�x?�ht+�}J��(�*���89^>4oî���]��E7úܽ���t�a��� �O�<�_&Ѓ^sh <�|N*nZ�R�7K�>nb�8п/��l	躥��i�`/$���v�>]������ˉ���M#�`|���0cm�8$��FZ�^��=�5����T����px3�����p+�-�%��+b7$�E4�N�i��jq��c�7�S"۷�C9
Xk���sA���0W��x??���{ �2�x�[��vӘ���y$ʣ��Yݙ�D_~�cr��`�$rOx��� ����	�6;Bٶޑ��ڬ�B�ܠ�	"�'���=���a���|�:7Ul�OU��f�8�����N�3���s'�GQd
g��xqտ:<�vi�w7�WT�{��yt/���V�p��r<J��cf��Pw/�B�.��eV
����L�
{M�p��~��b�H�yV�M�̩SQ��.�TP�e^Xdr���_��@��G��	���v�t�ֽ�G��L�6�T�
��"�va��T�����L���m��aQ�f�B����'��Ɗ�V�l��%6���=��Ɠ�{�l������u
� �|	�t&����?#bW�������˻�Ӽ�`�O"J�e�p8�70���U{��qjѫ�����la��e( ��"^+I!=����J�\h4<0�`y\L�a7���+��[b�?[q�Y�/��3�Ga���n
�P[˞��Fڊ,o
�R��]��hD
hiWNO�x�vcDA"f=���)�9�j���;s�8 �� =�Pg:�26��#��e��ʜj�XJw���y27�5�.�-���+�o%8��S�2LbHH���@�Jee��iqP�_�s�\��	&e~���Mi��f���n~�XOL���<b)�e@W:��]k�NS��������Z�l�Dp'UK�`����^Em�i"�E��}���`�?��!����Qo��V}7:�'Ko�������d��_� ��^d�=�I`��������T@N�I�pУ@�֙��S�Zqs�o/�!}��Zd�X��?����p�O>c8�Ţ��j�l�u1�3O2�~�1�g��]d��+�N[��de{h�z��4�@���CK4�y��0���]��e�w�$G;oR6�i�4���j�s���o��^|���k��o��c�{A����}�-� ��5Y� f��3�y1�lWn0I�)ܤ�2���)�ӃG�D�WإF���]9X��h�$>0/�GZ�C��~Z�0��.��=`{M)h�3q1'��R�T d�\z�h�����=�D+ֻ�tDzDVC:�����Ql�j�8	�Q��,㐮�.W��������Q�V�deX1\#���D��y�R���"ˎ�A1�EBCI���I��Z��1vʗ��ǂ���1����J�{aCԲcK���8&&�hh >����TA�ad������Ieo�T2R����� �t��f%Z���W�јp��_�U;�� U&�dme�o� �mЇd���ӦuP�SЫe��\?�ɺ5K�ѭ
���#q�o��_iL�����W��	���9&n8s�.��,��Q<>ς��,��E�A�h'�N�g��ۢ|�'���J�ǧp(��&�V�Í�ad���s��vU ُm��^ژ������j����	Ȋ+,N�p�$���I*�/�<��t�	ʗY�};��� �$�b���&~!���vb�
�i��_ 4�t\������,�rv:?�� ������'{<a�z}j�s�*Տ��{�k�_�;u�f|u������p�b{đӥ�'���W-)���.�
�̦ų�v��1AP<7��4�(���j{��9������ۙ����t���ho��)�S���V��1�A��\��y��P� �դ�V�b~�nʋ���;}Q��.U6]�`ut����>-�1�ڪX5h�G����(�O�U6i��d�+�:*�F�.vCJk�o;��ީ9�Ǣ���D���#��K'֨��QR��÷�h�,6�[s�5YE�^��=�W�L��p�Hxo-�n"��� ��xX��Y��e�کr'׉t�XY�fוH-5�R�bN��(d��2�RO��h�D��#%f�B�4U�_O6�L��LM������?<��>��d'a��������h.D��lN9vh"9���.�q"��"C3�����Ǳ�U�F"����U}[���u�/y��O�.��~���>0��߿.5�Ț�N9����gʂ��]-����-v8�����7[ތ�i`�<�[Ctn+�X��E4�����@8������h<K��tՈ�+�i��L��V4�t�V��������di�SW�Й1�ޔxg�6���r�s�v�-|Z�	�6��s���h��'x:6�(#� OM��Yp�P)'2`��.I�a�ƞ��R�ujp�%�S�����,��v`<�j�U���D���u�]YW菇!�eс�\a�k��� �Bh��ֳ����qǖ}��!���B<`�V��W�=L�)R���ǅ������r5���*��wc֮�F,�4E��`�*����ϤT���	����W�շ�rW�׽�e�����F1�#=�\q4�&�~z~��C/5��!\6M�����
R'=>��H��n
}�����`���3,��ӊ.UM��Z���o7W.��[���dw-���׼J���v	�F����Z�К���A�A'�+�al͎��Md�QB����]�̷{�\Y�����C_Ӂ�Ik�o�lX���ҭ��e�8��0��
��tUܰ�;p�pI�)e��|ޝ��06Q�u�E7q�JǛ:�U�|/ns]9g���՛.Fr��;���K�F�BW����$�%Ǟﳜ���0h���on{F���-Rŉl~Q���E�J�b�at�[J����W�9�#Yك@	�A�8c�.I&��m	l�+�T\��@��]�����#>Qc������"/���P�W�������LT��<[A���`�(��N,�'	�l�� ��t�|f �'A��3�ׂ���� -�2��u%���K���R�������ڜww�����s̎���8P�_�b%a`>����%�1N����W����X�ڽI^ъ2�<8<"��jF�3<���w��	�RbUFv �qC/�"6?�i.-Qݘ؛d���8�i�� (V�K��t��uq��#7�oi$���@MP��f<�JfNq��
Dzv�<�@G���K!�H[ɦW��'�C)�	�×M�N:(���U�	��ҍr����r�禯W9/� �6�5��T�FP3�Tu~ҾB�ł-�sVy}�w���ض��u�Y`���O�B��	��r3�p`I9�(+x��EK���U�j[sQqP~�k�L3�j�5�x6=6�_H���ätw�L�Cþ��k�*�^��+�����o�E^��鞮K��g�:�g��j��n�J���1A�k$TƍR���������tW��>q�\��81
�:�\�r�cl��W�)�Ȏ<��N,�V�p��6�M��~|H�:�5'[�0���:�FٚL*$_�4Y	������ש�'�*��x���1�X����O��0�nq�MV���q���K���f[.Eou�i�#�f���C\��w��7rs�|��Ų��rw
�5����C�5=�~>+ˌ��;d3qC�~	V|Wt���G�(�|
3ɛ8mQ�2V\~���ʺ�⺄����������θ����d�����V���/�%��E6,�����g�|��8�%L�dNE�9�w�83w�|��`��������#�8�g��*���bCLEb��ð�z�!�Ѫ㈃�t*v4���%1f��v���
hR!�!F�P�7��>� oD8l����
�-�Ԫ�����
(!�ĺ�=2Y�cN�f��3�l����?�]%i�e|�4=`�k�R>�Vq����2�PW�e}�#𠚼��^~�a�@�<��Ytp!�Vf�e�7S�@�5}���ӵ/�" ?��A���.4%$	�!��[BCz#��W��ݘa.����+������ja�
��Ŭ]�ٯ�L�l^>~&�Յ�j�b��g(y�E��1R-|8d��\R������wl�Ěx妬���<��ʿ���#����,��!��lf�r�RF�`Mxlkԛ�n4y)��9��� T��v���~ݗ�������oL�!�33T�4�(���H_���LڭL�-���M�p8�m��"���`�'kA�N3�]-"���\D�6�e�wg�aGPT��I��ܗƑȂߛg�XN~���ו܊ۣR?�����:!䪋�ٔ��go�����1�g�Q�r�V-�	eL����څ�qfFPTX�[�z�[~�pRh� �K�`���tn���?�̺��� �l赼g��}���n_x4�<�<��<%)E	n�'A��Q��?��&�֦͑��P�%��i+�8������doW�y��y�ٰ�b�?�d�`�!%f����F�]EM���+�F��m��EX����	��u�f�����,M/�tG�'G c���G�v��� f����f�Fi��Y�(�=G���'[`�.NC]�8��u�uB�馈��)D�>��֚e�L�w�b�(�?F�"�̓,�X;�Q��sF�nJ��~�V��@��e�F|C6Ԧ�KY�v��|Lgʍ���� A)��#�w�����E'�n(a}}�L���uz�w�rr��}{8�6�!�[T���W�.!�����e����`�"%άP��Z|�2K	������D4����N9��r��s��f�Bg!�L!�,#���?Z��4t��o%�i���s&˰�K)�lv|��	��_tz����J<L����O��M���+��.B��������|�ȁ���Nm�Y~�28=��^�QjW1�ʹ�-��$��}@�Qg��7�<�E������+˷X�������}xs�&9F�q���|'��Gԩ�:��{~�m/�pR�%=�v�d�Ln�|�L2�S��]g!E/`d��tm5:I#OJ����얱�����ÔH�2eYGӦ�H���Z)����t�!�pƓ���G(+u_��=͆Ƭ�3<Ud�Iɓ����8������~W�qÑ���ķ �N�<�(�k��|>L�O���$⭥!�T�2��H�sq�Ts���h̵� ������s�3�����J�07�ఀf%�l��2w�G�6��=���:1B�m�a&e�򍅚vZ��W�ZW���L]���y�P�ͦR����i@��kJt���NN�S�4l���_���*h$NO��t���g&�j�����:&t0X�kI��_���֩��\��^���#:�������Pb�����d������,�tz����="�w0e����4[�	���ο�� aA3� ����͑�~k�\�|�����x���έ�E?�������Zxi�8|#���A8uVk1L�[J�롊��򐴸��Kc�8�m읯��h�����<YI�����(�� F�1�h@�=G�i����f�vBU���4Z�%g�Ϲ�]������˴��� 7�?�sS���Zw��O4T�?�)��7w[uȼs�BiS��~���� �v��Āձ��G:����N�b�y���(��n7n �y�(8���|�s/�)�/�=`)P��5I��#F��$�)�E��)C�&�˗�	���o⹔�h 3:���wx���|E�e�*��{�E�/�#1ˑl��ŬjK��!�D�"�䌂v^�v�皯����z"�ˢ&�ԇ�*C�1P:�kQN�ffFw2�Q>���E)�Y��	����$��5�e���Y�k��Sߝײ��o)��}��P�f�(�-gM{�ϼF�b��_s<�r[>����]��@,iLd�~����w+#a�-�*q�Sk�R�O�H��o�#*.K-|"1�λm3�,�G��K1t" =�@n<0��D6��� �Z�k?f�5����[/��<�u\ye�O24L|����'�i �W���%�Z���m�
n��1�+ҡ��k��+�H/W`a�9nJ�������褎�4/v�-d0������5s���"Ԙ�<�D~�&C��ZD��\��+[�-6���q��r��e]����o�0��6�����!a��1^dn�&�T3�?_�.��E>Ɍ��]�l�0c�I�5����x��8�3���N�����Wf��L捌67u�_4�]a�}Lɲ�g?��>5t^9b b��>g`7b�t��g��`wl���q�?��&��ޑ �Qǿ_i>�3/܅��@�uǑ��j�/�v�����RQ����3�#����nz������k�A�/��올`";�_V�B�U�st�j�j݅�A�\�> ���pVs���m|��%�lvY�#�Tfˡ��d��:�P��g�'4ט��>�8��h�u���9�G��j��
�Ŧk�1|��V\�S��׳� �ZC]0-Ft^�ozy���-�G�UA}��PdI&N�����"��*<�<4�G
9��\ 
�5�C�C@��6*_��4�%PGڔ9JG'M�*or�:�-��xa󌈃���-������U����⎏5��.UMN����nѕH��sC$��UO&e\�a�����>����Wy`<S�֥;��~�Ǌ�T�%� ȁ�'���b5�yC�acUO�>��IP��o�\5�3pg��9���a|1�H7(�W!"?I}>����0�is�S���b�\I��,�+���7��"�? �5�� ��n�&}�A�j[�.�8D#���=>�A'�9�����кhȘ��H�_\���>��ӽ����s�}A��[�������(i+䘌�(���G�=T�$��߼$�ChI���`�(l��CS��X��@Ҧ�{�iu�_%F-@�W�A�=Qǧ�~��Mx�:ۛ����6G}�0���ΐ�]��W�0K���MqfT/Le���'k��.>���C����cW_�.8�7z���;���0reoJ`DJ��'���#ꪔ�\᭗��]ٯ)�߽��ێQ)�X�k����������|Ֆ��1�UU���=�W����5�@�ci5qs�����:����R)�ݦp(��Pk�8�"�����i�bYߤ����T�hG�,C/@��</�Z�?Q���3�D0v��;!������
��K��4�v�	����[�|F@�K��su��ý$��2��H?7p��ދiF�A������2�8C5(ψ���DjrfzE}%�&+Q��*��=N*§~b�o��:X���}�g��L�=a�:�.!��%�菽+児>K��FoٌÉd��{���o&�*�"�l��a���
	_�*��m%��+�a�|hޫ��b���}u�Tʠ�o��֚��uxa�cg���Ǡ��JM�ύ��B'9�!P��5����.w� D�2�A�3��$�yE��w�LV�����y/9i�4�,Z�Q���"l)��{Z�B�`��!ɧָ���>��!��#�	��'���t�E��W�b��V�׺�?��vd���N�iWZ3Y�m�Vh*oP��Vᗯ��V$g�=6���Jk08N<Q���&wULDc8���$-1W"��&ku��� `9���<��'/�VƗ����$+��*�|X��E�;2�!�S@�ܧ����t��⽗أs�1��Q��{�p��~y疻�K��8�=���,8*�.���՝��K�P�g�:$:�0J���;y�{��m){�d,�9F�
N׎�U�}l��X�,J�I"��bX�����Q��{��׏�d��bA?ŏmֈRmO�	u��Ȧ��U����*�0N�.z���I�E����c��;X��M.KV�N��i��g�
�iyW^�XH�_�;\Tˠ��eɧ6,.�93���!b}��i���<�S3V����q��DQ��F����$��/��cF��$�ع�.֯�'�cJp��^��ޠ��C'���|ӌ��ۮ&�r�nxL���oB�ɘ
�m��� ��O��m�1�=M�8q^��3���~�>��ao�&38,@3���$WW�sj� � �.m8��I�sFPw$&�E�3��;@e�yϹǂuDg?�n������9��b�r
�s�tqY`���|��O�$.����X��u��[�@�=��14����d,[o��IlRa��SH�M'��c������;��(�\�AGra�H�8*�*�zU͹�t1���A`�!���M���8���k���-¶��?Ͻ$�G��I�.@��V{E���f�-s�>�x���+}���YWԂ12���9���|p�,�����>S�H�ҵ:�
��������@�(�zz��>$"��t�K�г�Y�5�N����	7�":���c�| N���DHkƑV���Hp<Ș ���u�"a=rV':DF����2�e�3�����:FX]ƹe����+a#�m4�n|'t'{|��DR���dux�'�Q'K�����Hzq��c�F�q�����Ԭ��H�_��?����p�3��KΉ4URR�J��E�T
�����d�����M����M�y������a��W_�gۀ�+�������sS�������%���B{܄�Y���l�M)P��	���A����\��j����J�C�Izu���o�ڬ��?��%=�k��~��ئbK��I�8�d(IQ��/R�6� ������U�W���	2ղ
w�`��89'��x"�៭��JV�<=�����sgcn5��%��v8\ޘ�mǽ��k0�9�2���Rtʘeh~�D.�=?E���]C,���S=�t��%6,�O�T�Y���|���"�A��\����u:*�_ݡ��Ƥ�uc�Λ&1D��Рx��A�����Q�%����7����U/��孑#l�l�e��z�M����}a1O!�Fa.�������^�Nk�M��p��^����%���ֿ�";�׵[��+L�2��
F#�<n�N�$��� �桓c��\0Ы�5kO��,U�6�v9�����W�Bbw���𪁁����kvֳ���՞	�8�����6����7d�`��hut��ql��A��zY\	��;ɢ�<CV�I�������I-�zlJ{5�s������lSVfoh�� �v�Đ�6}hK�f�����1�~��@L�2I�:�r�e��3'@�e�`���竑7��4�!�u�h>e�sqhi!�4��������F�T������"�E`b�3H=Ydb+x��::�yw�cm�MB��qͷ���TRԉ��a��Ţ��Bi�pһ�5X %Aܼ����'��>�Rp>�Ai�7?2�3�WT�Js��kg0��J�9c��i���#Ћ�S�`�ϴ��<gH�{�f<��Bg�bp���Vf�M�n�2Z�0S�˰?�mϐ��U
5��W��$/D�Z��	�9に�6",����5K'��ZĊ�a6�E!6��1� 1�)�Wr]gf�'̌�����R�G��Ԙ���w�K�	H�]l�0�c������˷L:�gP<E��U������$V �T��=-��|�����	�`*	*��^FyY�߻��"v��ӵ-Fn�0�`��[�ڨJrt3.B~�Z���9���YC�(�]���[�{����Z�"��	c������x��{A�DJ�C����Wv'a�PaI,�v�F�w�g�ER8 S�c� ��*}o_�G	�!�WEoH�uOH하�2DC�&v���^���
�kZu
�~��R.+��=3�ޚ��7��w�
�+7a,b��������Z{�.���xՋW��K�3��Z�9�����m���c��z�b�w���g�c����
��˜FZ�R�:�(���"�zGt�_�I�+���:A��B
`4�"��Rܢ�/ ��*�s2�kb@���s^��C�Ϊ��P��O�k��H�Ae_�9T�W����ȿOI	�C����߽H�GҌ���5�%��UW�K3��lD�ԾL�1���5!�������δ���28��e�N1�x�}�!�r��?�x]?.��f���+A�p��;��~	s���R��)�r�����㨟�VT���;&�ۈB�d k/�9X`$f"[�oۖwX�#')��:'S� 4-��|F�������!s+L�{Sа����]�2u@���x�uw��/c�g����~��k�0����ā�+����4�e��� T�IV�a=1`�P���9��P,��s�u��f�;���([��:M���\j����8Kr�a���`5���m
�;�L2�h�����q�0�YQ�J/��?~S���n�k�ʘ'2�5�Q���\��펴e��*��W��ب�u2��B�q��%k�/6!]�|�x��,֗��-�u��b�����Z8��4���ګ���g]�	F�%������7h*Ah�ȼ@ ���7n鹱����"���몠���O��S��1ۺݷ�<�$�'vF �^WA���:h^�ǔ ��Mls(�2�9[p�ne7	����J:���~���vG��:��8w!��`7��[�U�.s�o�ψ��/V��7��b�[xU#a3�9|��* No�b�݅��'���H��&qEYh�Z������,89Y�%9��G)��� �ӆ�F�)}G(�}9���M�U��l�?��)�YD��Gc΢[��!��t$�ywLEZj��K�
��<|��f�
G�=�������8���T�.�7��=ֲ�&P�i����gK犲�||�
S����3�ˑ<hĀ�чDD�p?�Ȃ�T�����V���5����t'�����5���ڨ'��[S�s&����<{Q��AhQw���	��TŰ��;[/��~�Dp�\1�b�j����/\+�y�Q����]H�kY�����0�$O[k��4���td�L�E!u���d�R�y葓\���������` ����Zx��x����I.��8��S4|��
@�x~�{U:< v?�_�k�EsN���C�L4}�%ჳ��*���v���C�Y8��bs�V��.f�YY�l},�p2�}a�R�\<�3��y5]	����Zt�޳�� �������:���K%bcG��%��$+z1@;#Z���c� ]�;  mʦ�=��S�ןl�6�E� �H:lSDZ�'�Y�t��"�dr�Nq�����a�uƎO�,�c�R�XR�P8�A�2�0���q�j�x�\�����$;w�/�@���B,܇FoQl��G{+�C�������q7��d�78մ~|�Nϛ�2^lr;Y��?���O�z�x�����ͷ����0�9M�B�5[K}j����O���2y�;��j^���68��1���n� ��d���a�u�����س�/��M�ż���wZ|+���"����%"�P�#<�Q�K;)6�ތ�z2\����FG�_��c������ϑ��I��$����|���=����eO�\Cؚ��(e���Bp���/Lx�j- ו������U��(��"���	���=��r��0L��]�X��Id N�Լ�H rͱ6�\9��6�O���b7hzu���m��"�⣍���*���e�����f�Z]���Ջ�QvO��sF�MF�f$b��v�0��5�T��Ó-eB}=h�k�=��}S�ܛ�Y��q]-��SAH�-�!I��i� A�����������Z"p�뒹�W�dh�R�e{FX�5�az.�_⊘��A��:6�k��Qլ��w��ݻ����	��I�+���h�Ѐ%��ޠ���郢�^r�<����yfI>d|OT��H�&k�9����^��f��~7��v>�����|�ívvF�i;�N�FUn��Z`�*h�q:�W���{�bYnm�7�3�������!:<�˰��/�	o�%�Z�w�#!���s�ï��8�j.�4��֞�hj�E߈���ij߯���)�H��6b������Ns1K6{D�@�8C���a,��e����|�MW!#K�����3����:ьP
�ҭ��>D5����J�z��Ĝ�5~W��t�~����� �F�K��l�NJ�mV^��
o�⺸���@��Ex�V}��#���Q��B�������w�~% ��F��"���O�:��GB�6��7���U�m���T�5A���<����|�Z��+?��;{���U[@�bɇ95��Ý;�>����4rUē}��0�Ң��6�9���|���1I�fz����:_OA_n�7C�ڱuR�$��P!�]�s�5j�����|����\G���u�k;��ymA&�K�E�i��7)���Ȫ�TC�;&��Ӓ�f�����XMߠ\��m��\ϕY�r!s�'�2լ'�'xw���N/���t���GJD���}	R�CMAF����kU�����X�����K�u��|���{]iaa��t���UJe37l1�W��X����ۈ���F:\���S�9���JA���Or�W�Tw������"���Y=���9ev����.y(���'�#�B$��MU���RK�,؁WrJ2���1� 
�q�כ)�|)D쿟�ū}6��b��A���\��\��D�{�e9>�a�j��:�B2ɌLxU�B	u��OG�~�lbk����nt�y��K@f�RbE���#�N3�jl'���R��;~�:P�, �ĥ���;�r�c�ς�&p��N�BS�Q��_��!��U%�6�/X�^��c���L��Wu0�������������^W���&
�R�e��e��8��s�8�ۖ��+Bz����s�} j�x��I-�Bs�.w}^���&������1p�=p�It}�,�x�(_��%����#)�PU=��]�O�7��=��������8���Io�O���Y����G��)�f��mS�.�]�$!QR雕�buRҶ
��2�>CP7�nVlH�۪�$rHoe@Ջr�'��ѕ��:9L���~q�,��Ay�4}�G~��r�@���d,�\XE{Z��qjڃ(�Ssq_�⼻w�qdX5�sH��Dl��۴�Ա���~���IV�=�vr����h��uWY b�|W	:�, �G�uR��%��	{=���SF������nu]vy��l?i�-)����s檺:\i��_��]���z��H���� �|�ܢ�ѕ���y�~�U�F9�s0���.�$/��%JÂ��ΎQ�@p�p�1Q8�$�i�����J��6�^��u��#z�p��
�L�5sǧì�fɥ�'>q����M���bH@(>מ��'���(���Dw�^VN��;a�p�mt�ީw��Ck�+u.Xj	��P��*��eU_��Y�%��g����`��QÛ�h�߬��W�;��:�u�x gjl�g���7c�(�٪nN9�+�TA8a�η��0�{���7����=�a���Ǩ��R��������:&q=�{��,)���o�Y�z��U@�,��݅ S��lS�ҶM��Z��Vq�ޠu��"G�E=Bz�/�g"��ݜ(�C�=��a �w��8�`8gZRߒ����׃�d���{�-S,l&K턽�S|�V����>�>h�i/rR������i#p���t��M�nƒ�*}�u���D���t}6	��#^�B��F�I�VV�3a�)ꚓl�-����0�}����ˢ;��ټ�I��MdnsQ"�ׅ�q�����^��]�� ��R�(�[�|�Ҫ}��a����Eݨ��,Ҿ O��l[>-�_��R��q �̱�`,��G"Z�OQ%^���74W�Q�����#�pT�<T�S��n\)�W-�.x���J�n�=������{`E�%ƕ'ce~j�_<�̖랱�I���5�n�O$ �
Fk8�v)љ��ž@*�p��^��ѫf��1���UL�k�3���ױ���&�EO������߰K��������`��+�ϭ��.aosٌ�\2MX�\��n}#.�Խk��,hF���a�>A�� ����%�߁K��l�����[!�U_��(T�/�N��i����T�rVilᘱ��Ty��Όq��^����4�e�d��Y��ӟ;�x�x�qV0o[ט߶��?̜X!u��Ǫ}I��xo�,G�JX�M������Bն&�:�58�Ңz8����Kk>�'�8�4iGR@ږk�� 6u�ZX�{$m�T��Y��ӕM*�Sm:�PXN2C�O���Y��!0R�g��-BX,"m��'Ĺ����-\��.�`��:�P�ڢkae6VaӸ7|6/��I\�N��4M�|K>���#����\�8���?�3}t���(����X�4��|�x��l�q���<���� ������� 2_�S���aܰ�?y�i��b�HW�$�]��s"z&�n7�-�/���Nr%!&, ��!����Ƞ���Q�9��?��穵5���`����������3���krJ�gӈ��}+����6�h�	��*�}OZ�vu�8�Khef�۽�o�SmI�LZ�4�Iǻ0MO"����%��b,���ǘ����B�j�s�Պ��Գ�#$O��\Tx�Qe�x�5�	����N���ȥ�
�44��(���U�b��;�>aS<�t��j��(n��kE�l�ʇ���N�؏�rn��{������k�yP9�sI�|D<�Z�E���OoH���|�P�^z�2W�)�e����4��]*�����ĤA���z[叙���䆍`�	ASZF%�̡�'ai� 3�TZ���������`�p�1��e�_
�l(�A�� O�R�T�lUX����ww%�T���1��*7��v��ʥ��Fiʵ؝���ݺ^/T�Q����� Ϧ�.�N(b��U��UE���'vS:?�������գ��k�J<Lj����iu0<�d�W�`�1!�76�u
�U�Bk刍���ʄ 0�C)JH�	W-�`�ܚ�}禛�s�0�g�� ᢵ�O5�Cd�Zr�,�[G F��o�4A�Ϧ�L�X�W؞��o�)�N�e������>���C5$�S��=�C��T�\�����$���� !��n%���͈�NR�����9uJ�l/�6%n��r �CXJ��A~��9�K@5n�z���T+�s}0�5yFh��w�bKi�Ӵ2����ɨRL�5�1�8��_J:t)���탮����F����`0���b����-���6�s��z���t�;*H(����[w����DZ�;��^Zv�*��Q.��
����#0��{�:���3G/��ʹ�r��"�ބSd{M�ߦ��+� �d�]��%�
q�b��������y<�ڄ��?����������G7�IC^����3�E���VN�m�Yk��n�a��p�N�'T
�le�: ���'���ԧ��k�]e<8Ƅ�b�Q�iq-?<:+畏L�ңzh�.���n]1ݑ�!��	D3���`����`�C,0����Z�*y�A�ƭ�j��H��֖��Y�ɧE4N �H���������Fq�����7�z7n��@���{�@Q�c*��9P�����r�
X�r8��)9�+�2��32��E���@�7W�$���O�0E퀝�)�'���#GS���P8� .�xR������k2����
OY��-������;���4G1a߇B"E5S7u�-Z�-m�t����{��%�*S��~�	I����Hۡ�1��ޜ|:�3�R4�Wu8NF4Le�
st�����(cɿ����Q�@(��2�v����c�g��n4'��Z�P�_��RXhQ8�^Ѐm�2oW]y,���g���҂|v�K,.�3"�a�A��݋��r��'�%�O}���N;)9���_�C �)�/0������[�}��,s��� y��!��#Nqnc���p�4�UIDWlA��ŀ�s�������!}��b�l��3#D?[�Ί���4��|���/\�/��B�ݥ���;��ɘ����-P%�^���n�gN��S�Ǖ��Kf��&��eT3�b(���|��R�#Q.�t��T�^��E�;�,�J����F,Vz�]�8C6.X�I��������]��(�Cb~֗�A�쟳TDe���=�q��F򧪊 x���B�v��/A��;�|ߞU�*�¹i���M.d�I:H�yB�L	�#��V��Z��ݓTS0�
v��BA )�;�8�����z���ӫ_v�1G��	�O�4�3&�X�R��"mcg�^��+V^�j����F�/�PϾB��L�����$�Kkl�� Ə�����u��4Ӕ��
�+�{6�{(3*2A�	y1��u �ˤ���"���O^R�h�N=Br�$�����]�QY�;��I��EǰTg-̖T|�`)�C�^[u����K�2!�<꯳��.�Z�Kc���
6��:="��d�XX�{����2Z���ߴ�I�5�v����p?�����L�ƥYoK:�H�j��|�����>�=�^C�̑���n��	jƇ�e����rqa�����",J�.�ܬV��
;�^%�04����I���G�nbi�3��b�����\���:�n�b���#Q�W��b!��,}�(�J�5�C�Nl7B���~���4<�)mde�&��QP�ZM���6�C��v�l����o>�ε�h<o�!�> XȽi�s �o����&n����^x�r��k ������ƶ����Go����SaKE���>&ބ�����ﵘP1�tH�ܵ�z�0oi���G^SaR_�-v@��Ȋ����y���<���S���烯DIjr'#}T��5��@��V����{��mQ<!��/v�K*��߃�}��]��+�0`��
��k[[9��@Z�9�\���s}o�
��ej+Q�����d�w[M*/�Z�!�9�T���7�������5�0����ٳ��{��~aN�p�������p��{��R�$3�L�f�<�h��Tq���*G�����4Q�G��`E�)�����nOKYÖ5N�����o�H�0!y��0D����Ј�`:��^�%x�7+<]P��3�8%ɨ���64��^33�e�>نᤄ�e'm�cx�y����J�u�+% w�r��&�]:������v��?L�4xA�Hѓk�g/�fSU��M��6�\��Ɠ�*)ds��"��|�0X#���)B�}p4<W���X;}�,3p�f�q�^��=w�z������2�7�2���d/-ԶkD��T:wHÐɏ�d���l�.A)��wÚ���V]����P\j�p����瑼�3���=�/He�+fU!�Xa��
Ԩ~W/�/�]7_!�������y�`B�u�aua틡�N������r�P@h	�h�aT*�w���aI��$:U����c*%�Uâ��0~��z���=�7mb�ܨ�2@����hT�td$��&������T�n�7x��A�<�ȝ�,��G{�[�#��k'o�{�P��1��!���+������2�b��Ok}�K᥷5�@��SZ#zQ�@tCd�@�G0&��� ����=7�S�F@��kA�XK�u��z�1�m�M,�br�6��I4{a�]GJ�v�2����,�|	9�ūҴ|���κ�=p��X�k�sNlI�o�0��$��@�9��@�`��>�]�Y���G*�3�R�QEP(9-Z{��_����O�CyH}��^���Z�,��z�9B�9���m�\��*�(DKVT�9��ջ�+�3#/"�,y�R9������qJ,�ѭ���|��F@A�&�O�ƨ�&���$���:���,�=�.9D
yJ��/�,������^����19�G�������L�{�d�� ��!���T��t�VORO|�g��2��Ϳ��e'�qȳ
��
���Z`I�.�5���A�Ӡ���;�|�t����	���i���(Ce��<-�{�z�r\���$3L����Fl�F̀E�e��5X���fc1�)B<s���%�.c��An �2����칩Z� W��XiS5�ΖNgq�c�M�&���zc�n�} V����{��]��!�����Q6�����U�\L@-�$����8饠����]!5t�YXp��IC�2�K�y��|��+O��jp�3<p�p�֎���N�2�z�$�0�/��s�Bg}쥣M������k_�u[�z,|ơ �����Ƽ�8cGU��DzK>)},��U�.럕b�5	�Ϳ��A�܋*?�����A1��&tsA7�ep?�A)s��^Y'�%d%�[�@���L�vs!���d�5��㎟��<[p�>�F� �R�cU�h�O�\C�St���ZS'SC"�5��u��$ď�Ӗ��$�/񩺕��ߗ���{S����5�}�;Qa￳�m��E�S�˸����C�i5A�);>�.��\_Q�
FA���"�_qr3F���U���4�t_7��CO�K��v\:�a8N�X=��W�cg����HZ��>�K�Us��8�OM#
��MKmeŚ.%�A}r�ܡ9������� iK� �1��Tpka��)w�Ҡ�e��� `�y%���MA��.�m�o��Ց-Ľvj��ځ���u�����<<8�烬IO'S\�J&�{��n�5�����%H�ד�����ә�:l3��R����e�Y������edP�Ldf�3�(�`������.�����k���ݘ'y�\Z����&Fv�ЈV,{��h]��7:(rEsoΈcu��'�^��%�H�~�ZA��Ʈ۽��=��Φ�*�/"hÅ��C(n�V�[01;�H�����4�	�)�[Xr1+N��Ƚ�K3.��Cwը��{���uDt �Sٯ�-�+��&۱�o��.�V;<�\�_كDd����@7���G�ZW�L/��NR?�_5�V6�3]/�'�N���<�����F�G��fcR���Z�j������P�ۂ���$4�fp��D��>h��T�=��yB$�� X<X�%�z�sL?|���0�}]��z��v�M�I����P7�]#@ye��r�P�8���Y�m��hT��RS�Ƹ��\R(**`}J�/�!���<�]Ĕ)� L���P�lh��i�ҫ�t���(��Ⱦ��1J��v���l3��G�ܵH�?p���0�M� ��1}������*bS�ށ �I�-Iz#��bo�J��cW���u�җ���9*�_i� ��]�J��Oۆ���={����k1��6)���ב&Y�``[�$���C����a/,�sib��7�!��`e���BAM9ȭ�K*T4��R`�΃�U�N�?��elp���n�k�e+�̦�O�$�p0{`U�������R��=zetbol
0/����5f�E�ɖ�k�I��Wq�������U�lN�L'k*�� �{ZI/�ƈ_W���Zv�Fߚ�E��]���N�����&�}�	�7��#�3��J!��-IK^pKO�L��BcֵT��Y��	��0����Nl�����[�/�K&fG�+S�����g�/�A�����{�J�#�&����
J,z��C�\�8U2���_o[aW)��}1��d%ߗD�i�P��ـ3��$�D! p�0.y��/E�����IK�ؓ"�[铼�P$��ԇ��/6����ѤۙE��&ĝY�T~�;�7y6��q&������ܞF�&�������}5:P�wڲ����Z���%ܶ\�T8W TNn���a�	��Se�����H\g�����O?�t�D(���FJ�G�y:��L�0Ң^���u�G�m�C�4��.Cc�u�{l��Uzj��냐\ti �k�1��T�f^]C���#荤}}l� g�YeqN�S�km'я�F;'_���Ip*q.�Ƨ>:��[���qL:�>�$���}i�*�[�� ��J
"S��
�1��WW�3��aq�E����-�Ly�uz�����	0�ŕ�P��%�-

?O�?�������Ƚ�@�b#8;�%^nA^�����ۮ���2�/�E�c�1��;O:�u�(��O�cYF���GM�[�����m����k�B�(a�G7��*AS�z}я�.�Fo�C@~���P���O�lPp������߂/���0Ug��u�=��j��2��1�_�N�+�h��ZI0�^@n�.�F�����e�+EZ��y��6����M`�l�2��o�ʃ�@į�8�߷�GK�d���Ӈ�V��X�؅��uw��qh���R%�0�n!�d����G�D~3�$Y"�ޣ����x�9�'&���P����Ȣ`9�А�
hz��fmJ�c6G�
>BL��0�P���j5�<��7'����2c0�^C5PR;�=������,�!�EU��D�=3���۰�7.Jr�9:��1bj�,b�~�ި���^)�y��ȜsnF�F���'��H��{'����:6$�x�E[$cE��|���QU5
�����S�0�u�-`}�֏k�z���+�M.dF��n$/W��8z���v'�!�$�O~{���=�qbբ�L���ɾɂ2�R����딚jX����W���8r�(Kz�?�hH�o�r��|�a�ܼ�/�3�Q��r���L8���xy�TV��hBt��]2
�3?�G�R�}�W���\��c���QBB��_�CϢ(Oa�o�
�;�T�g��:�<�GB�MYWթc:�L�z�����meYzs�ס���(ĕ�1��m+��8IWג���;��HK�6�P���G�A���Ļ���F�&~VYSOd�I�R^�/��&"	)�*��y�H���
Ac���^�	o�G�(,W��(9Hⲙ�����onK���[DJ�DdE�NQT9�o�}���с���z$��J���}�B./x�wc��Te�,�I�x}�A�����ltɕ���(fFX®�6?@����b۞Q<��P�a�P/�u -����4�13��d|�ֽ��J�ة����$�hN��o&zD�>���~\��a���{�r��@\��w1 �H��Ι���ď1��
��ưuk���m��9<�6���4`�
�-������y��pa���V���8��,(]9���������~o����1\�KRH��HDG1F'��Z5�t�Y�\����5{������=���;2���`_j(ܤ���{R�k��d���Zբ��H
��l�zA�/�݂�q7�c[���^W��H6��R�q�7|��(,��| �w����(vE��b�����-%M�넔�^���Տ�H���x�7(�)�����|m�韵EYZ��R�!�6�&���^����@���
��i����Ŗ��D��
�4��,��m�^.�"��UR��8�v�9v�0)P#h����<
t����a�����q��y��@R�fM�#��v.b��g�K����AQ(k�%vT<��dVOV@(�z���d�QYWg��w��O�rv�q��C�����ł��P���ۦ�����f��y��ɐf�Cn;��5���є�n�|(s����i��𛾡�㘁�O�hb�h�$�?�|����a��b�Y�����㒽���g����{>�HR�֭�eO�&�7\�����4j�4ƘL:���E�L���o5�	E:��ẓh/�ˏH[�؎� �.
��{��Ԅ���a��V�4��x|�� t¯q�Cݓ��r$�]y�<a<c{j����z��B��V��~k[=����~�#��v�H�7�
!R-�k�h֍Ik���+W� w%˷��)�ٔn����M�����
Y�>d��ް,j/b ���#	�E�up�!g�*w]{������k�$)��� ��-8Hm��-
=�&-1�b�r{�:u�kfZށʑd���ٞ٬TG���<c@=��(�G^�D�=�gl�R<���@��p���Z�6I%��ǚ���hePEz���	�Q�O������Ɂ&�Rg�킹��� �g�ެ]�^b�NV57�ʊ�.L�e��*dV�0�6�݋�&ɁF]~�ţG���8���|��?�MnF��z�X�Oi^�/["z��:j���f7�Eū3fD��4/}O�fJܩ=RlP쟻t{�<�[8H��T�j��Z��ʆH� �M]��#@3��Հ�Ԗ�!�܏�DC�$�^U�5�#p��&9I������Rځ-�<Ӧ��0"�P�\��oy��Q��$@��k�s��a�/GJ��Ư�k��^@^����o�+��k���~�on��A'��a�3;����Y����"5���Dc�Ů4��N3�D�k�t���=Ms�i�)��S����,����<b�-�4_���I]��i��NsX٧V����@)U�.��5��;XS�..��fVԛm3	Cm�j�U�WN��F+D%��M�pe�ai0�����eQBk���F'�l��?�����a����aWCZz_��q���;�����vV5ځ�p�g�N�"�(��s7�6	Wju͈L�Ir2-b���z/���e)��$�b��R�I��9�3_z2��T�8zT������i�n~x~]lpk�!��-�-�v2!��Ip�-���!�T+�o�]_I�C5��-=��/�� ��Մt9�kV�z(^W�:�kJ3 �G�֔Y�aSɵO�F�.��.�������d�"����/��Z�0S��[MA��2.JH,,���&��z6j#�4HG�+ݨ�y�ˆ7��(2$G��Y�{\oqHY��
_�[YlF�G�O}F^���B�F�L��y���jŰW�v��<�Z/JQG���#3�Y1g<�F&�yIpe�l����3�`T��`$��Ŷ���se4�mJ¦^_�����>��� ����}�X(!bJ���($H�ѝ>��:�q}�rBĢBb�qX��y��h���5#�,�&��D��������!QH��3���%�i־�ʹ݆�*�򸭼H�cY�'x~|�/g8���6����}f)|>�e�����U��,�Q�WO��eB�B�eb�
	����?�ԧx_��=����;�x1Z�s��{·.����N�<�m����F#�!4a�ɵ���)0�E�&o�c�%��E��hY�p*�Q⁚9H�/;�Q�&�r�dC5,��(��~�럎#o F�"�����d�|��٩ *򺪇�@�9q;�^���mX�㻫�r�ؗ/!�;����P\vR]��oԌ�g�n��'��=g~�]��P�Z���kZ��$@�s��o��~����˂c�D�J
x@I�a�Ij�nPԍ� �(2t����ߵ{z��O��pHe��j����,Z�=tz}f�+&�	���@k�wv� b�:W����'T��3�]����3��:@~p
�Y.�����6�Q���A�ƦQV���*(�e,������[�b��*�f��#���ZϙձQ��<�e���	��N��j%S��cV$"ѯ�40:�m�O6{�NM������5~//�獇�EV�B�^38�*T��Ҋ�����͉�������+�`���d<�u>҈` ՙ1�uw�ꌼ���X�I��(l��T� ����ɔ���%��XT�vu�����췿�J�fL�N��Y�|	�@*�w~xNG��/��f6⮼Ŭ!:�K0��̫�ɢRY��j�=�	Wu��^,#��?�W��^��0��+1�:ԎAԁ�.C��R1������+H`m������>�$������q�&�U�hRK�-��� �.SPŮd9�/���vBm�Q�e�t})��nߟ4�k��|�C1����`�K�oEP��������(���'Ѓٳ�hƤ�E�Ǵ-�ї���XK�͢�ԃ�ƚ��I����GL��]���tJL9��ol����Oa�m"�|�Dp�֙���|DQ6z�
J`�{=�Ms�>|%��0����I4��V�k�n�x˅��#+�Va��+�-��<���~��#���@�ń)Tk i�Ma^Y��.-�i�C{ͽ�@*MP�so�Kv;�k���6�N�s��X W1N��Ƃo�g\�B���;*��2fǪ��Ǘ��ZLqR�� �k��K�k�D�+��%`�vT��L�9:D83(�����E�R���s�e�=�S��0|���T�ҥZ����gzAY���n9MO�"n14��x���D�pZ+�]��w�s���o�����/��5������b�H>=���|���.���[i{]Pj�d_2���8��`.�Ih�TP��Dsɿ⛄d�f r<{�ζ6^|\o_̬y�Fn+h�g��ʥ:����<n?�Ѹf�a���>U��l/u��-��W���+ɾ�O ݓ����f�q
��V�b�p��eRA�-�H��PA�MFC�Y��M֖��R^�=b�tA�����&���+���͐����s�7.�猡�<��g�Nmu���4���i{F�1�m�$���+.��fؠ���|�(��	Hn�_A����MY��R��7F�ss��A��NP�G�a��_�nGY��f]�?"���[�� !i\��e�.tK��eq�-��gʨ.�y�ƮO���Մ����3����]5}_>� jþ�Y�VVF��#�iV�������Gn��/B�ܭ�^�@B���o�}-��\��������υ᪸1�l�ƍOhtI@�v[^��+���+i�c`K��C���[�	��Cl��R}�Ǔ!mU�!"7�1�B�z��ۘ��|uG�@'u�^%�{:��N�H�I�uf�0독�\�3�CߴDxX-���5uOx��oPd���D�o���/��^��.Ӎ���+�E�AY/)}0vė����pa'uO��p@���D<b��yG�HVg{�Q������l�37m���ð�j,�U�ʇ'	�:����W1af�� �F��2'ͥ����$��V���u#7] �]H�"v�e�m��
����ۅ�i���ͬ�C M̛z�A�PԒ����8�l�~�}P?h��Gr����3�]ᓪ�zH�^�&�y}�b��؇��9�`Dlc2+��}P��>*H$:_n�zvkX��GO�]���áa1ޣ& 0j�l�rI;
a)v�t��&~NM)���n7X!o8�îi��8.�Qٞ䲿�l憒�1��>`E�������-������)<�,�c��x���q��8�,��=�2��),�(��0;�Kщ�aO��Ӝn��n�:�n�"��Կ+a�x�����2����w:S��o��&H�gk�"9��8`}i�1��d��ک�s�}y�Y���G��H/-^����5C��T&�'�?����)�_�#�ƬQ���P�VF�VCn��b��U����׶/5���q2�);��cX�>D�]���kG��J/�����J���x��25�|~��k �w��Wpg]B+�\�(��Y�v'���~����-�wZ��..C��F8'����L)��m`��X�)v?��i4���f��O�v��6ٔ���-��g��2����'�o$r�1��{4	��ݤiuL��|A�"��]����#�k��I�H������Y+K�D��T��au6�u7vۓtO��l���.Rc��ݝ5�� /�2�U�d�dBf	+��i[��Q����t�P��^�����qio�_BJa-���V�4�wC��w�� ���ȋ�B�Մ�y��t
�Fb�1�鸅�����^���j��!{�A&U�
"�����)H��ƫ�hg7>���^Y��р�M���F7�����Xn�>�|z,`Fo�H��%o����Gc��o̔����H���p�2߻�;��0���.⸲��˜܉;�Ǎ[)^%��I�2�
�I
�܈�e���fj�ԣ:���YBO�B�����hCmxܔOY�
"��s��,N��&���ǻ��D�L�!;�ٛd}��Ց9��oLЂQX���}�?6�Cr��Ji�UG��.z�����\��Y��?��f��~�9���ߏP6ϺX���}u�b�g�h���j��M6��X�㵱z���}�'~N�8��(R�p?j�(���z�"�2��%�.�;�ɣ]b�=h�Q���1,�s� �׊�^K�)���J	%��U�:/UIR`���I"oc%^)��#t�:��.��|�"}�D��\ᮡ��? t��%Sر-�jW+�CXa�~0eKY8��$���w�U��������ʄߖ��)Ma�y��G�����щcH?��g�'��켿�a��5CFD$e��\�o��ag�O���@u +�$s.�jh��Wd&b=��~>������s�$�ӄQ�L�wy
��WA�L{�R���}E��9.Q��V����=V��.��w��P4�}�4o���:�	��Y��ݰm��Umٟin�-��4�����n����=xV��M��V�����^�\��I��@V4/��PW���O�����T���P�@��
w>揌��d��%�E��}Ȏr�������Z<���3b������(;Q4�[�:�cQ+.�n{}H�A�nVs��"�T�;y���*;��vdd�vq�e
�Q{Ģ7���c7qGb
�bs��˂��(���Դ��kQK�)1�U Ǉ�I�Z�C0{u�ߏB}&,�[77��Њ*���E�G�G�fw�F��0�¼�sZ�'�H�q��C�1-������,���B��Z��^�-�tK�Z6�� �h$ad� ����F�]s�4�&���0@�g�e&��M�	��M�+Y�PF�?erRBK�`�|&�@R�r�	��X2�$)J_�o���O|�щ�Xq�$�<�z�	�ߡ�{��6@h���;�TJ碹�1����.�VbpM�2�]���Հ
?X	P�uK�ɍ3{3�{���/��;�K|#QY�U����e2���3��w`�R�(�]6��\eH��*�F?�V��\9�0^J�S�:Pp�"{���s�6������"&@N�Biʊ�M�����,�r_��P�>�X6}27�b�4����n�2��Q|'����.��Nɮv�(P�L�ÓX��H�C�	!n�/�9��<���:E.k�[�uɖ�ݱT�&nA6��y�M�⫩�zR`���k=ںX�݇�;A�!�׌t�<O�P(���5���R�ѳ�le�q=W��Ht��h� a��5=�H2e�f@��I'���?i�b�̌>LsHU�!_��h���n���a�ٰݍ�7�-�B�;v�)��@�/��Cx7��6��M�c2��?�6�~����ʢG����t9]:��:�O�Ԏ��D���K�yл��65�w,�ƥ��.:��o��t�Pz�m>x�C�+�{h��^!8�5����@R�erU ^��1|G+
s�A(d�Ԗ׎����=��6�7I�)0(��*WУ�&�N��6dS@i��C-"���AAůw�_��)!��z���|h��o^y�>�~�́���F����@m������N�C|ۅB����һe`NY�d�{F\��qD�A�i�y�0�1�{�MId��9���n�B��$赌�,����>n��x�Z��az~���k3E�{Lt���s	Xd��C�bv�} ��Lى�@�[皱�{`#��Î�L~iN�y�fÐ����d\d SckI�����Md�R��r���6�����}��h�UXHg&��b£�bYׂZL	R.eYX���ȉ�
9�%��dGo��e��Œ{랬��i|���4��_>��YRr�b_�"C7m���\q�>�r�&��wU����m ��>"��i��2�H�ݰf)�e^�	e��	V���.s1:\��e"�G�GR���'űG7$m����*#�u*֩�� �- �@'	��G�rB���������d�%Z�c3���Y���'��j�(��	qw���@��Q�i[�B���h*s���<Ii�AD"�ۢ0�jMh����C�(�%�dLdc@���r��$Q�C�'(�'�(�u��Y�ב7V$�PX%ͣ�nmj�#��f��<����S6HÀҿG�H��<Ic�v-��xU�NB5Ev-����\#A��XCe��e�5�ŻD
�b�����lICwu���œy1���3�s��%�vѹ��B�*8ޗYp"
���K��5��$'����je���INU"En�$6T��@.�Bo(���A���y#�������}3�e������2tk��*��^���F�G�H.�bcb_���Ӂ)��pof(����[�X�k�:�X�ЈPo��Xy���lY�������N���e[Y�����9N7�!\@A�F����sؖ���#h�,(�;W�7\,��9����:���_�j?M)OFN�N5�Ed��1e]��\��#�����ZS@�����+\���O�J\6BOJ�v5lB� ��K�Fi�J��$�N�HE¡��ޓ��X2+�eEb&>Ҙl:��ed���`��o�Z��D?_��6G�@�r�A�8����~v�0#����������X
������9>�������皴�Yʓ�*B��p���xc��;a�y�����
Ԭ���$�����N��䁢=���Q�:��<W������)�2C�?�C׹�o����^ee[]�D'ޅ��HU١���ar��p���t �=�p'�J,����}��d*�J��!@�Qw$�t|����\aS/��t��p�Y�?:BUl�5�I���PM`:�鹇��(Q���9�k�&~(�X��G�1��8D7!�Ml+7I�܆bJ����px*�'sVKv�2��p��Y0P����{��$i��Oǟ���$hs��9F�L��u?��t��d�O됃)r7�J��Ȯ�W�SU���&�Gs=��q��f�ƺd�Y��m����޻*�5C�v]�뜏��\��)<0������������ڗ��Xo�%���^<\�Q�8�e�u��D�S'��dd�r?���p����(��� j9�����+�Q��9>Y����3��ЊyA��K�?!<�+s�p�� ���zl6�F�'��г7�,Ź��p�'�v�0��菊b���H��;>g�|�9��^l���9/���3�3N)���jIu�a���C�V�1��^�k����D��v�'�w�q&��~sc���T(�4��5B6��o���O�@������y��v)gDx�E��>�IQ��$���"<�Hɳ�� u�4]�� $\{j��y�(�g�{syiS�X``���r�:��k��ژ�0���l�Y��5��`��[bh���N���HHx �����Lp%��)�I���9+j�}��[��(���� I������5u�bA|]�E��#��Ca��\��[�,)�W�"�e�V�I�q	���6��(A��qBr]�<M�?HLOV�|�t���4R���̈}��O�tw���f��$/�9e�q��ΜF�/ �!�1GD�錎��97���p�O�i�)�Z�$-��VOHDL:zK��|�5�5���[���ԕ^W�5�	�e�>�X�S��aq��tM�-�x�׭_Kr�ٕW�����[1�u�ⴏ�	�ճMMʝx�_�C��⤜I���b�oՍ攡,�,z�l��,��\R�����2�Չ��B�2���oy����J�C��]�����$���#��4�j���]��y3=aՃ	C��h��[��������à��e���%0"�`3'	3����G����-���*r)�-\5���$�=�grKr�j��E���?-k>����y)gR���_�'=�C=����sؤD݇�.�5VN\I��x4F�Z�|��3��5e�P" �m�-�U�ʿ��-�����KE��ZrNUIY{Rbo2ߤ�틇-��o>|Ҹ�����n��>�K��w6��8�:~p6��R�o4���GN8��P���,�2�p"GhZ�8}>������0��Z��9���⸅=�����ҽ���3XU�'s���^<�?�L"�z7��.�^�ė�,t"��s���B����;�J��+�tR�&0��oj������#�bP*�oCBi��]��\���M=�ZM������
�<�T	S�G�RL����,B�D�:an��~p�,|�~7w��k����끑BbSN'�1J#������o��H�=a^Gbi�_�6�{5Cyà����ܰߛ}o^H�4e߸�P��R/����WU��z�\Uê&͋\��^_��IN��5��&��XT�2g����@PB|$fI��'nw�f$Q
%Tµ� �1~�����CL=�l{����柦���y��`�O%�P���\�|��:c�C�,V��>�u��㇡6&*��:7@)�bb�;�Ϫ�fn��养�9M�*��'v�jR��5����}�B�-:�n�q������ �o���\{oF�&^�)8�_~�qbi��Y|С� ��9�Օb�v�ݾ�������ECMI�ӥ���/���'ю�黀.ލ��L����r��om���96맬��@��!��6���z�)�p����Ls_���%%5�1q�Q�(��8L��۳@~�`�������?����n��SM�)����焛xȩg�% ����oD!�<�3��8�ψUY�8o�eZ����ږ�M�C���(�mjl�s]ۂz��fFzk&0���wX�齪Ẇ�W�K��+a�E��� d3��7�׍$N�j�׾Ʊ��>Gو�%��o|`J��#�+��5��o86�\9oS�Qg4_��'�����84L;�����ЎМ83e�������3*cP�U�2��s�t�$���.�.T� �CP��"�5���E9��ن�9�xS]�̞���BJ����yFF4�ݦ���ٍ�8ta�y�kJ}ax$?�Qf.���4�Cds3���T㡥�-���dN��8��Þ��c|�WkAsp��2�è�v�< �&�|�Ɇ��.�P��r����x�񕎝@��b�t�l������旺�=~��.�$ ̶�{g)��g�Z#��G&���'�7t`H�Mi����Hn�9xYd�.g�J�*�㵳'kP�#�b"�Sz�&$s�&9��IS�9��z�
/�+���׭�|�=�\p����cD� �����~�Dc� T���"~HV�7ϫE	����`�%�Kc���!q(h��JPƇ�w�H#����"'̤�}mYr}��9F*`��h�>K�zWƷkw�F����1��Љ�t�����#+$��8 �i=���U=��K�'�-`��B�
׳x�r�]1�G*c�иe=յd
x�����M�W���%�#6�>�o�΀�c�<�}��=!n/`W��PW���� ��\Ô;Me���Ȑ�9�!�5����?�	$Zoa��������մ���%��;�ȱ�y����l�v�{�<㥨�*��z̖������Ę�6Z�9�yzW|�.γ�#iE�&m��^y��/Ox$N���O�F�nZ�݂M�%N��m��������RMF�~�5��Z��=��p�뼄1W[��Yq��3�f����@��S�%�&��co��/h�~i+�c�)�b�Nd$~���_���s�Y��"�0���o�*ڜǮ��X)0T�ޱ�3d�4�>P�R"3�6Nk?1�ZΠ1��|���9��r����Q q��%��H'4q`��IDM�X�[ڇ����	�m�`�����kљ��^1���]��q@�Lb�F��k_9�b�����n��kp��0�	�5Q�r�M1ohI��k���9c	���O�
�j��S�bo�]O��.J	``ݎ�;	��T~��&�9��4���lS���R�3,>�1D-�=��Bݓ��Jo�(�!��\�VGO	=�V�E�}����e%��p$�3t�D>N��G���BJ�T�K�#�^�*Ju<z��������
��"���	���W��Djv������,�u��w	��������a�a�c���>��I�I}���V1�dL]I	�A��q3-z_��?�&43a�Z�kQ��ќ&��b�3�=�lN��a�U[[&=�,��\�S}=M�����EdK�p�*~�4�Fp�4�	�!G�EEv�N�w�R�G�2o�֐�G�����~�p�Sn��,egPGk}%pv"*�V�'�Щp��o�V�=Eʮ�R����,,�`�0;퉡���g|4����bX4Z2̃)�q�W��<�o ��N�����N��Zf��Ʊ4�]�T-����OOrcPFϲ���[�E�?�Cy���4����o:1���k��@�^���r4���va��+�w�X�д�"ȕ�\߲lL���6k䝯�<��(e�xʓ{W~M�θ���,�*��+�`R�J
���o��*��2��ZQV$�F®�m'Ƈ����s��h�g�W-��(����.q����B�?K����
ș/Lמ9׶��P����+�$��d���
k7��qx�\�`w'�(�]<ک���'�T��)�^�V�"�}
���u�X5Xq)<�R{�G�=~G,���Zmo&z:d
�1�^��D�[�E�}H�%U�ꚑ|�1B��#0��L�N+R�o�鴫Qw��}�N|#yێ�Ϋ�}�i� g3���쮺F8��+�s6h��z��H;�]5�Y�g�o<��}L��I�Z(!l�qa�{�\��0A=}+�Z�W�|�ԐRc�M:���za�Ek��-/��F�]{�S�fX���Q�u�t'�T�菌y=[�#.K\�)�,	O��meNLΏF�t�ݭ 6SRC��aA���������)�����1֣2|󎳔E`����Vd��-U]� ���;��7*֓����~l�Z<"@3i���O��m�D/��QقX�汢��S~��tK�)6��VN/�b���U^U:�U��(��!�vUf��WN �3���hPȠ�Ic�Y����=�Sʋ��i�p.o|v=�+�YD��h1��'���N8��U�N�c�G�T�$�ӛ�Yq�.@�TC�X{��Sb��_2P!w9՟�|��!�!'}M�_<�c��*��d�DΊ�*�ǟ�>�Yz�Z�y�1>~���u 5��e���������)��/ƉS���F�sJbD4wK�[iB���5�
�ݡ�/S��)���8�����x�6\�2(�r�N�5�h���b��,��ܮ��HX���j�������h̑�s��xlD��A~�U��<�唋��1�_#P\��׊J���O�
�ʳZ$�#��*/�!��M�"y��5��N^�a�B 'X�\e�@Wp�� Fj-fQ8���J�K��/�f�ht}&��B�O�{Nf|79̝%HB�&�B�����xo���W�?¯�����LF��v2о/,Xh�5f�6�䴸�t}a�}` ���'����]�F`�&e%.�"A79�Wߍvp�j�9���ϩ΂��2Ȼ�>e!�]4�4��#m`z�k�B34����'u9��?�*x��3Gؕ��]��vc%���T�u:��쏼�Ƣ��N�I���	��XX�����J���S�x��M��� )2�����Ɇ^r��$�@d x\���@�ߠ�|����^qPh7C�S-m�x��e�x �>D�R��N|I������US��sM�b�eًC��c�6����.;f��?	�e�/�I�u��W@7_�d0�nR�����t�6_�sT�N	�hmVߜ�S��*h{��hׅ{��>�+�wSyJ20��_����k$
��t
�UQ�0���(2l92����D=�Q�9���<�=;m��iB��<V���}z�5��<xJ�[��������u���A�v���OHԇK�G���'���	���,F�`V��o�2�s�tsK"X\6i���uX��k�8ki����6抑8����2,r��ǩ�M�1-�����@BF��6ZT�a���������Usi^�r֟�)�Gc��h�P~M��9�|E�G.��#�L�q|�9R�[H���7 �,5a:��A�T�鶡�|8�a��\ C6���/1�i��6ۃ2�]��K�Šd�֩�J�:�9PY�u�&�a�����d'��/���1g$��ۃ���Y���0jն�T!���z��RČ�v�Y�R�л%����Ҡ�
A��d*��U�L�px]��5-��&���A� WY�f���ȧTA��L�'j����w�?V��`�n�C����S*#Aa�,uh��w�*�|��_v9g��*W����j[�F}h��g;[�rӝ�d����<��)��|�H;�ֲueZ��"jb��C�oK�l�@i���r�1렫$�Y>�R�ovƿ�$�>6�Fٳ��7��ٺ��*��a")��&��B�����M����1U
��<&��;�9�:ְ����<�ٺ�~�e�3����Y�<l�����=y�\�Dqt(V�>G�V���?�R$nYq��zW=���]��[8���}�>v��(� �DŅE\I�Հ�V�4Y&!�����Y XX�ؤE��Gq�^ ��|��6/�k��^v$#f(�����/�͙����+�{��h��!�0�����X[��Ś��#��J�e�m���c<�P�_='��	@u����`:Ե�����xRHڪ��澜zx�U�n��x���6't*d��8i2����7z.iW(�3o�Wn0�*�EN��d�*�(ܿ�"��fF��;���u��cSf"����N [��yHJq#-���[8)��Lw2��a(t#�?��D�]T���d?�>�_-&�l�2�F}ƴ�S�߲c%��?:-�{&�t�Y�Sg�P�s���8��H�k�+���Q�oWH�(�\
�XR{�$$(�
C\�j��\�ن'���u����63��h�&gSbr�IW4B
lJrY��N�K>i��gt���:��涞mw��d�~Ʉ]�O(m#@xmh���C�V8�ϊ/pgH����R��#����A'��܏�D\���5,���^`�M���O�����$[G|��lm��K��O��@mR{�x����Օ7�y)"��="dq8�"M�J������+-�Y�Z�g��
d^��
Bղ$�=��ej�XH��U�4����6jX�U-��pjYw���!R��5r�P�$��S��� 4��D���4�k�	/4y�=�-���UrE��}#�0p�WL�gv�*��h(���k*�f;{��.�/��u�]�+v�>➜?K��yk�� -���[#�r �c��������
�>�r��=m»�[�;�|�9��t�����	�SO�M����ѵ�;9H ��E?i^���?eIz������#�)y�1���j�ƥy��&���3Ga���?�|m�̇[�GM��Vѱgn�����8����� 	<���?��R�)}D5��	���Q�C��� ��Bu2�H����>���71*|�N�G�b�!/�{��bօ���~�+�uʠ�f�MHyc�k��{	s��� ���@��׍%7��*ɜ���P{�!_�4�kkH"�7}��ح��H:���y��CЮ��m�څ���Y��+��5u�������_{η���w���5]Bc�XgE��Ӎ���a{���rǆ�3�Y�o�WT6|�z/��GhZG�V�6<�
�U��̽ˇ+����'�Pk"��!����+��)��nBVb��D�C�?��r�h�}ԇ&���ۚd!�~M?4����%Ů�����s9��ѧE�K�	B��x�N��=���S�f���ڛ^����#H��ɷ�	�(왬k�����L�$*���Ќv��Nq���Xip�/��e�Ք5.�(R��a���5}��v��y?�Ĵ���.Bc�R/A�^PXj�W���2����I��"M�"��hbf�o��9���|ԁ�:�wf��D�'�|�񰔅Uy��E3
[N��;q4�d�[ ��c���|�}��u~����!�H6t����<�V�w^�Qv�[wY��"fΓ5��E�G���B�_��,�E�$������@�v:���"#�q�2N��$�����i��0.(tR�nS�{m-����hr4�v���X����_6�0����%.T�Mkc?���?���E�)m��ƓX� o3�����VH�[�Q�����+�w6eQ-]�*q��q'I�lQ��@^�N�4�2�<ݬ��@���h�@��q���Ӈ��B�g�o��ܢO}xo��50�un_��Z����{ر��L�&y���ǋ-$?W$��²�JJ_2Ms0��<���a�W���|�Ȇ��Z�-�Ao�t�T��䗯�ׁQ?L��M
��W=[%�u�}x�K1��]�"��IٹBڹ���{�*idO�qMPAJ��؜cҏA?��?ů�C* ������%��TXtt�8�ԏ��2�?�Q}���S��}[�f��q^J@�{H�4ɑ$^�9�����je�~_>nڧ��Y+����?aDF�:��m]�����o�Y����{KזXF7>����%��;����W�mc�c�d*"��[��=�LdD���+p������^��L��K�=K��C�u�ʜE�0��bH����Z�fR�19C�s`Sg�SK-�
��%��q��@΢4
|GX%��`�j�"�y�2�����c�T�&"h9���9���/b )F���e��L���>�m`V�RK�N�l}Xd�v�r�< �W����:~Pz�Z}�A�ju�5g��GN�h�A�x�M6-���)��G+D���U3I�ê&$Q��;ו�#a;N�']�E%�-O��_JA�.�?� K�S���K�F^"���M���D�^��|m���2�ۅ���MS��Q�6
�b�o��n�B��ߙ��7@tyT�R/��7��!ξ,z��ݶ�/�Ծ��E(��o�����{����s�h����V�Z���R8^�x�W�ɜ�!*�lx�����j�F�W;�T������xM!O�@W��r2-vK&�U���貶b�D�V�j �E���D:�,$�A�����	g������^�OS�]͸� �6���1�����6e�k'-^�S��]�j�����'$E�%�$����ފ3��9���N@~��G粊��#�ޠ���Zj�k_!�{SYx�!����O_�^w{+)�YYM����ݯ̱���aE!.�ȣ��9cc>��3K����Iw"-`lW,��pY�@@�]D$��D"�T~@bD\P:X|h����w�K�����t���(�69ؖ�w���%�߿:/��8z6A��NaLus�VN�R@M&@��L��Jg�F�i�Ep�HA2YW!���� ��1�̒0��hl3��m@�ηy���9�N5[ea��y������`�ҝ:5�B�]�Ċ������@n�]�;�r��2մ��o�c�KO�"��|�����O�/U��(0�-�������^�'��g����ʘ/��f�ߔ_]��Y
�Q>�kRO��s��eP��"<���c!qBi�gw���������%�� i��u���ޜ�;����u�Ԥ+g�sZ���.���Ё��v�gp��eO�-,��]*�����[!��)�V��t��K�w(�c=>�!'�v���]P�`�b���n��@����N��X��
��獺a�&UW8��r��i�Z	�qj/�4��7;:��7�`��2ҧ)f[*0	]��T�A6����/��\���l�B�[tA��c;)-b��QY�R(����\Q)O:n:�{��Cjۋ	:~e5]:�G��_~��mC��ICR�������;��aBI<�; ȶ�`��PvbgQ-_�]�݋b�oV p��Z�4��c��6��|������k�Q���B4���h��N���Qπ�)� !�Ҟ5�������ƻ�C4�\Ez��P%ەX�(s2�F�>6��"��$J�Xމۉ%x��{(�i��g`�mP;�NI�g-�i�o$/
j�"=e`���{�y�n����V�2�\�6s�.[���:;�m@��ҀLC�I{pk�� Kie$N��:��\��i�ޓ�fP3� �֦�MX*u7I�Y�<�7׷��"2�V)�0�+t+�
��cY��ҝU�Vń�[�!��uGB�h�t��=1ֹ�lj1#B��W<��؅�m"vY�6ۆF��+��f�;����?Й���A�ݡ8��K]��tGH�����1�Sg�&�:��F�����ʤ�Sd��'��݄˧���j�.��3�>�;p�{@�/,�巇`��΅�c�[#A+��B
�Q�x�����Z�"��@��P�a��b7��u�	��(K0�Ġ����ԙ�B�&��A
}8�k�٢#-���@��`c]��6E�J/;&�!����ᶷB�E�Q��4�r��x�/�ǘ�J�ciN�^p���-;]|t�jN�:�ir@ݮ�o��� wUIU��,}�[�4�B��� ���9�v~���{�E=~[�7њ��	���D	c���IΆ	�\���$s/�e**۰H�>�}RK_�"�e2c��/Aky]��+"�{� �q�2um���T~�@1O�$�.�c݇܋A����b�q��	i�^���0�~E����-#��M
a�rշ��'I�K����;�TMX�ŵ0ht�ڈ��	I&��B)��6l�0�3��/�"yG��ASY�S,�O�����8Y�t�#�0$G�%�o��Q�=�Q�.�᝔�줴����{��H�nN�=�������4X�0L��X ��_O����6��P��#3a;��jSy�6J	�*�Q8k��bY�3R��bS԰<AϭE���)�ӧ�<�c,'�Mc��v�4��<i|�$L^Ɖ?�;��ۛ��(��<�=��\S�$�Q�JXd����и�쐲X���Ggw^ĥ���z�l����i�d���/}D�w����
!�\��� ��\GZ]E@�߰>	�H2�x���u��Q��܎3	ZM<T|�S���2Ay�s�}<_���)KZ!l�,Mc�L/�X���ԋ����V������ڦ����[��zlG�.������x�;9~�	g���Y��E��d�u�a]w�&ez��z���@��	��)�nF�ї�#p�!��J$���=+���s�W:1�����ھl1����
X����n��`�*t�]�,P�ߗ�`aZ����)���Ǻ��A�_u ap�W(��I��;�c��!�pG�Xi�4Uv����1Lr�lM:Ns����Ǽ��(�=��8��� )�Z��nߢ7MM��4C�I��q����Z#��
�fAǞzG����yo
NY��۳��B:��InfG��3w�40�����5�b�����TJ�*���C9��iyy���!�1_e	��{�=�����3���쥮��3D=7�����Al8[?�X�
4�HRa��i46T�7c�w)�B=�Mg-o��Ն�Cau�]�Ɣ 
���N�;�
�{RoQ�%�O�� ������j�:;?^��2_a�㰇!��^�ܖ�,ZwЬ1��f��� |oR�7�l�l�]���֭�˗@�:�v>�R�Q����/T3aj�	^֙4=ԴD �(!-�=g�/��5��b���Ti���zZ �+��AL��~͈ݖ/R!�m�-��5�r�ͻq��('��	A����v9�Ot��J8�����/�z|"vG�Zn��,��7�Ҭt����K9κ^�⒍��
�7۝<edFǺ�*�r�&n���T/����]x���C�GSm��D�
}A�o�Zwx*��a�Q4� �K��B�ʈc"������T��V��L�(�ID�/U��-P>�2�m�QE��	�j��\<q�7<��N�6F�������<���8Ta���Բ[��]Rѩ�mҒM�@Rg�S5���c�\=�i��Ɇ`v8��d�s�q�m��k���0oQ��!�'���!�Y�y Ǖ�l��$������f�@1AuW4��99� ��ron��OQ�:��Ϝ��'A)Pg��
�\^����8HSn<CM���L*����3#Y@���0�΋���@�1$�`�
����d�G���DQ	�1������1�״�W4e� 4L�os�ew�Ѵe��z�;��	�~@!���-��ρ]H_!)�8s'��]f�V-r`ٿ�F�Py3���(}4	\���������j<�R)$y���Q+���;�|.f��s����S4��֍����a�WƱ��B�6�#���*��?}$f����yT*���H=]Z����teޑ�oO�Qb������_0�@���$M���//I}CR�T���c.��m��j=��	�� �Z��W��j �]�@�E����$�_ ��W����Bqn��T�b�i+�����J�n�_�&��\.v�$��	�j��Rаp?���8�{n�k�&����(�g]��6�42�hT�WA��o��ދ�Lp������z\mmw�l�����w�� �Pl�솱���A���'Q#1փ}"`�3�/�����-
	� 4�/�`��o�JW���~������O�i��>�C>�{D�p?i�z)��ю.N��O��hB9��L�_w$Y�_�#�	�����ي�"D��w��O���� ���1tkP���F��b G$)�)��V�'PM1Z�Вs�Z?s�+���`�iE� &1h�F�F~���������HA�"ǯhǎr��޻>�b>WJ'o��S�8M�bë5 ��$1�����2���S!�V6�y��e4�x�tr��VD�����dC]�k"��p��($U���[�|�*���ozz �������w^�X��4S^���K�ק�
>�|�c���z��р~���_����-L�?��/cԺ����1�@:��q�����E���l�F}=m��ǥ�Ɣ�9�G�~f����U�e��x-��3��X���X����ؙ�;�q��4"�z`ک�]�-������bgg��W!�� zz�5:#��Uw����ş�.W&;27�l���t��ȝ^�����p�=�joɠ���T����b�Z��m�{y��E�w�eN�ޏl�r�t'��B.R۾q+��╙����#�M�W |��H��"�=BL�9�c1���gf�`��u>��B}c��m�[����r�TI��	��C�v��$�y7���d������jO�Jޚ�SP�-�9�?�	�<8^���`#Eѵ?�n�?Yy�_V��>x�6�??=َG�!��U�
2��%8��3��ɒ�\�����P �ތ�[Q�tNp��7N�P� ��j��"}w*(�<o A�3��s���,�J���u��|^w(K�u@���~�$"<DH���V�kﴩu�$�_S]=�to�36q��
3hbu��9�C l���rV4�c� 0^���;�7�d���׹�]���:��|�J��WZqm�Pĕa�q��O߂q�ѶXC�Wd���}4�R5���:#���"���J�e:P�f�ɘ/���(���H�}83�����Z��똤��f�39
�'&f�g�}YD�bX ̈��[9�D��O?Qs��:�����$=+�ni>�iy���!��d��!KzD�e&�g.AP���M�ϯ�Ul���q���)�y���ڇ�f�C�?ƒ����R���R�B���r<a���Ui��fv�~u���۬�}Rn#�$J#�P�5�\�T�j�L�ު-�����j���2�=z�W���{O�֬EX(ZdM�����I�4��`��DR�Fo��#��%�y01۟�}�̙s��D��b ��`g�@܅T�R�dc&Z�xt�d��������s=�_�ߝ�n-��<�a�/�5�[�,^^7/P�e��|�]���>�j���xxJ�����{���Ŷ�4f���궣�ڙ{���cP��/���yZ�G��hч*��+|��v��˼��Mw���d�=��f�\�/���J6t�i|Y�'$��P=���"�g����X}?�1@�㴹�(��䣑j�֓�`����]�£�hU����L.L��\vVq�+�.Ѕ�M��v�8��@�� w�S���*H��Cb�S�Nnm�j�{�����׹�Қ����b;z/��Q�Z5��ŋ"y�[���g�q�t�\�c8W>����&l�H�=�=�`�#"Ղ�U�U�]pQFa��ا��"ȩ�x���A��].��	1R�6���Q���dD�Ѹ/���M61��)M_�ѣ0W�5	M�S	f��]���\�^�/&��(�c�(C}&;�x��&��A��X��O�|���E�_K
}�/�L�yL%-�6J��x����0?���c��LcC�w]�6���D_⁑3��q�@鐅�6]�
��?�����z0��v�cLv&���J��� ��+v`#��1�� ��	[�1H+#J���[b��&�w���JkK���V�T�|"�Y�;jf�2�O6��H�ݡ#m=�^�[~�g�ˬ�h/��8Z��;�P�,����_��m	�:��7��Z'Ee�z��A| ~�s��&�3��b�Tnz�k��nh�*��ԑb��'	�3�?�m��CY�� �!zO3��Kq�k-�
�_`ee-��r�O� K�b�����bqp�Cx�7��Ig!3�'��%ɂv�e��ϓ�]A8���;�C���Mgl�`6�H��?���A��� 	���hC8���Lt-���S�(a�N��P��>z{�(S����y͙]�^mG�"��V�.]�"�.�����f�8��H�9��$�[pkM!#)R��9�&����m�ߘ5H"��}�\����M��x����-���$4����bT���5زbs��k��m&��Z,B��!qu>��i�c ���2�`@{����;�}�a{��&�f�i}��eveD�>;��?п@�p����d�^_�d�<Dyȥ���Kb���	�ZQ#)hUoR2
�����C�����̳V|�����ϵ����@&3���(��T�h���5�95^U�����,�^���6vy�C}�� �� �j/nߢGi��s}K96�pO_�����h��	�NݣQu��Y7�� I��HV!;ݙ�G XE�I]d��L�M׌��9��|���N+����|$)1�w�%��Uk�=��rޏ2O4_H�l6`p�@�� �y���ԕ�N��'t1}�D%u5&^�*�q�Α���L�c�ml��Ydk�t?Nٌ��(	U�U�̞"v~򲆛��9�z�ˤZX��5��:Di2�!:GL���.��-I��
��Pe���5�" ��
�<�/t9�+�uӸz�u��B�� � x7� o���E�N�m���\`�z�Cd��uW�ŷ������s������R�.`%�&���w{�@6�Um3��N�q B��Ƶ>2�Z\��K��0���c���q�@�n��n�3�����v
�GbEa�}9̡� �!@hD�kN�s�S7�G��m��bb�����)FJ��?$Ű�Q6������A.�L��=�m�*P�ViN��ϥ��m�����q�����~��T=�m��7�ZkS_�1Ud�8r��|�eq�"��;O�<�AakM��>�tO'�rTݫ�%^���VX����V[$)��g_�t}{1 RW�GG1t��p>�߼�*XI��E�+���U�/��2�����x� �'�!FX"-��k�rɎG�r�xR��ɢ��^�e -U&F���:��Q&?A�$U��6Wg�dyrj'�1���~a]l:��g�0?���ڼ~���4.��L)Dx���+� 6zV=Ec��xw~��)�-"��nh�}Bf�5l�j��k��p|F���a��T��F��'O��Y���X�v�k�����}�<�/�J�H��>��������d��eM|�=�����;��3Cc1���">J�A�À��[�����m�1�x�ϼl������Am?�։���+u^�g�VH`A��n�!2"XÁ����%|_J ���ؤ��ҹ@ �q����썎	�f{�~ǻt���]Ex9KW�I��~�ZgL���ѝ�BeX���P� �^I�Ez�� y��A�ɏ�}P^eDS���kt�ɏS�Y*��B|���%��g�}!KA}��򿆫���	�j>�_t�|j�;��ӑ�4.�Y��=FBZ�hd�Ow8q��鑫����)���
��H0����?c7CW�A�Y$�ꌪy�7]�Mq0��<���;;�Q��V�"��)!W�w`�2��@��AV�(�g-�!Lt獞�\�c�+,Zz��ƙ\�[����K��C���ՑFAݥ��+�S꽭S,R*h|yQ}~�e΍��m�"�+�v��˼Ё�e��􋤪��k+S,l��ϥ"�����r�/xU,��5?|�kY��������_�1���^�y�Z_>��S�<I-��\��F��ӷ[4n��f�0a�%���������^%&#5�a�֋�*��c&�	�!T[OO�fh�gҞ�Z2�8:q4(�z`���@f،��h>P`Zwax���-m����sQH�320DA�C�nŚfM���ҷZ�3)߹�,Nꍡ
�~�꠮ɩh��BLK���'�-�q�18���̸ ף7UA����#���޷� >c��i���fq	7BGd���eV��H<r_�����`��w^ I=7��!��1��I�S���7�1�� E�e�,�6��fOI'�����ؓŨ�"1G@Cש�|��nz�O���3�<H,�v�����|�����.�%f�E�[2������4s�)�T���F4<�X�yx2��:�����(�0�LQ���e�£�����e�*������*��@��`���'�1_!)w���\~\���5�̄L���WG�4ϭ�d8��{��������t��@:���8���FM�g�+`z_TZcY㞒6��4A��s�`n��F;PQX�(�wR�{������7��12�����LI�0�m�\_�!��կ��r�o���Y�����h�~Тy��$
���c}�9����֗A`�������)y �5!����Y�(1W��0/�8qFR��ay��n|�=����*�a�U�1Yz8�l�zS>%B�hmO{_��1����5vP�"N����� �<
I�C��I-ڼ�z�F!_U|�I�N*MU��#�t����n�1phH	k��?e,)0i���o���ͬ@QK<�pA1�`&"�cv�����$X/�fi���(�^B���ө%I)9O�H.�`��y��ऱ~@�Jyy�_��uj�����QR���;��Q
q8U�JxUu�@<:	����ʫF��~��^F3��W�o�����^�N�_�����R�m"��o	�yA,�!��αu{m���I�}��>t�_;ok�f�|�ᘮ� fF�4`�ܶ��w�#q�>a��I�~�KcA|�Z�A8	�k���Driݽ��$r�4���״l�,�EŽ"	����Ye���X�,�ȷ�C�^���#�l}��'�L�A	�<>p�L�A3��������p�Ă�F�����6�s�@-jC���&�`M9{H�~?_Z�`Ӄ����P�?��6���H�ܓWMY�'�����t��ކ�LHѸm�����m뵾�zVi�C���L!|��|��wq�8����~:=^���X�I��$�$0hl��r�����t6��)��1dXa���������y�e��0��-	�Vb�UF�xhx �!h������?h���~X���oS���[pSq�����}�r�`��-	�,�/��@�Q�0������g��z9� �!Y�}�b���l8fW����y�0��s<Uʱ����ZO���Q����~����g!��ik���Am�Y�BR����9�XG��0h]?lVtT%�ϓ�Hd\R5�v1l�c��y
#�L9��Fӗ��	��m�Փ\��&l�����.]K��*%ҽ䈑p]���wgx������ȥMN���C�j�����	m�в�Q�t˝�.јfpk�+�A��,/�VWb�ӤT��چ)��_�C ����*6Bv��0ت��#���h)0
���V�M���V�\� mȾG
�W}
t�t��K�#�Ftu����U=;�|��b$��(x���h�M{��p�v
�c
�߄�L��܎OI��b�nB �x�������/�K<���'����ȍ�/�)lX�}�J��M�o*p�[Ы�P±t�Fjo��t~��Lݠ��c��P����g<�ģ�\����-ײ�aiJ�[�WC�b��i"AՌ�������¿�E,*�Vb��I���6���[�����&�/n������[\7A��P�^�Tv�6ew�)���h���^��z:�J��aG��Nfߚ�Цj��F^���zG��"՛�cD�a��#�D!�|&ŜV�r��,��3	0vJ�a9�0Ab,e#�&�&�(�UE8��%v�R��Y���]u ��Ӆ-�{�11����L��%�ob�
�c]�C�l�Z �mCs�M��^�pE�6���3 4���3=�x�����x��b�A�u���E���/R
M�� �^�n�+�N�>�?'�M�1��м�uT����x3��}[�{�1�N��6p0K��Tc��d$��N����n�|�M���3�̃�F��ġ`t����^[)=f$�Tҿ��H�A�[�b�{V(�+���>Atƣ���4��*7��s�&	�bJNh`N�����v����m͡gJ�i[  l�l��Fշ���s:0�XTa3\���RE�g8Ӌ{�Q�Y	��fU��VM�ƍ"fl�
�B��E������X�IZ�W�6\'iG[���|�W�]�̋��[C��[��l�1oTE�'V��i]I��#�b�g�ѝ�D�n��e8>�/�6vH��O�5s�����܍Ŭ̩�U���?����aC�v���^�U#�L�dۅ̌m�i��ea�Vu���9r��h�x2�C�\�?Cg/��G��u�[�m�mr������T接��?,�0�V�\ ��9�6G�i�Z�n�b� ���aaSqރD��Dh�s�Ğ�Lgh0��'qlym�:6�������K~{ʤ"��-���� N:�~��%ݦ��?����}N9/�u&�*X�V�f�/�Ro�N
��;�8D��X��X�b�:�G�"���/�hTF�$�{n�G�̡���N;�#b���I�@Ȏ�� 1<��m�O�&L��;+��L%)����Kd*C����n8y��Q_�迭Z�"DϜT�jh�铧,�v��}p����	�gߔ; ��rP��Z>79�?x��qݶO���=Fy��Y�: ���`����ˮqK�ܸ���T&�Ozɯ/S��u�M�"ʨ���JQ)�ssa��q��Dp��a1O�TA����4N�
m7o�8Ri�M#�o@�Ͱ���l00�b&f╺�G�4+bH�և�O�(���U�� �Yq�/��A!jJ�Qˏ ����
�
�=���{�"�ap��=3GGr��R�G�ސ:OG�hh��G~��`�p�*�rH�̕tq�_�l��������գn�����\kS�eT�Q�ȄƐ�X�*�S�*����#%kj߿��,{M���H����T"L�5���v��K�y�~�+�mȤ�yk�&�xI����aʡ<��N�R���9A�.�D���ޠH}C��)Eo�ߍ�l���������_��,�2�1Y&]S�'e���l�1FEb3v����8����#%�l�@d�@��H�����if?Ai�j����es�e�����H��w��{�g�E)�}B��/p�<D�܎yh������}��y<~�!��Z�*g�c��h�MӠ�5N�c�{���ѭ7��S�D:��Y��Vě_�@0�L���/+�_���Ł诓E�	����s��)�A���� L��AP⚠������*�iΙ��wO��
-�9rJ����ú�o�gj������[�����Y�Ud{�ɺ���-l��/���
p����zV�����>�������e�� ����d�����b�����![|�3�9S�@V��}����fD]+�A�8��ؑށ�m���L�C8�?x���`�0U�9{f���;I�+9̜.�T�E#+s�6#��gK*�A:�� f��A��~2����I�}G���lG���-TG���6S� ^8J�^�*��[��䳀��:������������.~�ֻz!���=)P*g���b}�^��o(��Flc[x�)�]U����?�X@���w�س��'Ԭ�?��9:�~b�b��s�oh����y�Q��ޝ�ǝiy18�%xG,��:S`ik�vd�Ip$�V�{�_*f%n[�a9i���Խ{(� Ĺ�.b�/����v�.�0-ו���0���-#K<+8�;�H$�ƌW���0�����x�^�c˾ޅ�q�{XؚL)~�Q��R���)��I���� ��ո5]�Xig���9��#���8�����T�_��0���r�����D�kL~�c|2��\\#�J���� �}B��o��R#�B��8P3�\"�����bA���|�Mm~C���\��������B���[�un���g���(�L��s�L�"Fe�K�I[h�>��+6����~QJ�l��ݽ.��Z��/a`+�5# ��f����9�x��t�[\P[�����'Cjto�4��ۚ`�MD��"�ů%8��"�*�(p�����2���=�GtABl�I�.$5w�5�|��}s	�cϝ{p�_	�I/��y=��;����O�<49�E���0Zig���*�f�CT��rbx��a7q��sqv*kV�xKynçZ��p�r�-�mq��F[THI�:%�W=�"x&ɫ�1�:�dV���n	G�]J	3=T���;!��E�4g�I
�����B�Og�9�H,���AdC�G��M+>e[��*̝���=��j�l�]�@�?��x-bA���^����t64�Lͅ�suߴ�����*�n-��ҋbR?9��� ´Y�#w��=0S�=W�.��8F�`���k�g5'mil��U�2��3�?Deo}��4?;x��k��a#�����E���`W]�Gvvy�\�8iTR!(q2�� d���_N�v*#��jր4���
��q���'T���r犣d�8���Ǹ�c�;q&���K��$��%���2���\6`p@��"�C�?n���^��vh�y�߯���	�� S#��Y6�GC�q��HtU(/��E�Ű�*D�q�c�X�������J�Os�z�q����u�r��/��	E�cϕ�S!

ӻ����N�s�CX��>#�O����i����<�@�m���<@L�>�E�s�!��-�%G�*]���
�%]�/��;[A�_R���IJ�XE�r�������7�~�)d93�'��0������5�=��
Uq�������^�OSnK�<K����z��v� B�`�{c���w��|ǫ��*`طw_I�Ͻ����B7
���`ƕL�����q/̄�z��B�� :ɂ�?�~�/ӝ�f��Q�è��	0{���w�җ�N���6�!:L����+1��XS���j$�	b�z�%� 3����!�E,����Z~
sC ��"�=��Jm�y 젛�ڛ�	N���_Dq�4,0|�;�A�h�2e�Y��2�����܁�R��.�*��S�[�Hh���\�I1u��py;B��J�1�j�����;�?�]�\?rE>
s��,�4 O�mWw�l�M�lJ����N�t[s9X"��<��'E�,�5��ұ�]ʹ������J��kᑉ�+¢��� I{N{j�\�`��6��As=N`���'y�8U��!/}$�D�s�pN������af��Rq8#������h X�A��U���[qk�Ӱ{�v�$�B����,�S�6�P�A��4�y
P�[���>�n��y���	��a�y9��>pu��n�[������Ac�,��x�n�+�G��=�����g�b��C��&�1����[�81Ù�_��>����6�R_N궜&��8T6�K�+Q��'Ãwh���ұ=�骂�[���Μ��a%Ak�[e4grAQ�t�'�̼1�����a��t޲7���U�}�+�����	l�i D�%}Ut�uSwI��
�"nZ޵ɩi�y`���{��o��bk�w0w��O77 ��a��W���T��&O���R�<��1�Ч���� ��9�N��_�	�v(�4
)���������܈d�f���v4N��zDI��q���!SJx_O��G��;\��EԘ/��\�3Hu)(�|I#+]v��?���L�3]��P�!���o�����{�������T�׊r�U �?�Η��B<�Ο�P]���ό<��Ω�K��OR��� ԅ�p���9�\v[H�F�l���5vB^IR��`,),�D���*�	C>�̅'9��U:��<�7@�eK�Qom��Q�BH�	;G v����`��=�B�N�~���O�Dv9m�]�n�5Tx������ȵ�g3���˪����'z��T���wm�Y)�(>��}�(��[oM��!�����pu	Mڌ9�B����G����֘*݉%M�ԝGԃ�&9,�H�L��c�`���^cf�x
C�4͘��5�CG�@�Z���V����ub7����yp*�7�����5�8���nݮ�?<�����2k��8��j*�r{2󗢁�F8��4��I#�����a,sX�+�p��~��7�l�R_�2źT���ni���z�a#J���&V�a�e�(�y���}�"%���_�v�`,�6)ٳ�Ŋe_wB]�xg+��NE��p��f�_%f*��vCd�cׂ�U�٪.�x���W�R=H4)�j���j{��붧u�3�%qڳ��՞��e���ٵ
o���r(<���P���� V�Z�����F����o� ��T���5U:U��ؓY<�XZ��5�y0�����}��!Wr[���/�b�9�W��I�����@��{�{���%my��->�������e�۫ ��0���IkM�q�Y��n��J��f����[�U�5�ޫ�
U��@5��6|u �QS�S��ړ�fJ�֡Jh���H��ߠơZ���5`�C���v��?�|3�	��"���^�ͪ<��˙?q�L��͌V���F�;e�Pʣj�9p�ȅp�ve��R?��������{6�b�O��~����~2n�oܿw�zU�EÚ������ɪ�)q���`�a&�͈`;1Ucq��t2�=��ق{ԉ�H8K%R�b�M�����Y�����A����s%�}t��S������U�c�z�9�8���W~)�V����
4C�U|�>�6E�(�2�{,&E���z݊YSФ"����E2X�����L�~*
Hy������F��e��Ce޹ɐD$1������!�T}��t>_X=zP�RZ֛7�`�*$Ҏc8'�R)#Zw�8õj������?�c�����JK뵝�%\�!#PEĐ�^�dɧ���&�|�+�k��K�?�Iz'��AĤx�������Q	2[G��x|.q�y��j��f�Xc��j2��M[�uz��I�	�d��RS{�v�p�2oDT�,�ro�k*�ϔÇ����Z+��&�m�V��I�>ldױbsڗ��ڞ@ ��A϶��wc��XzOqc�� �'�.o�"�����m��uq/�cy�-:�l�qā�#Qd"�K�=m.��l������FȓZ����֕`��#.�{M�$�sL<h�� �b��;>R�(6�պ4>��u�X�BT9�K�hR�'�H���J��ѵ��$�=Q�aP��� �pC���v��D�c�]$�Z��9a$�}=��\��q��K9Y4�����o5x�[7����`RS�,�Vw!d���y�(k�'lDm�:��Ǳ�:�{B��^���Br�Ӈ�BW�Arc���	g[�A�0�*�����݉��g�)V�q��Sp��7h#׬���kn簪E2�VlX58�[�̜���kH�&�vf��:����Lz/��uy�G���Q��A�'9,�Y~A�/"W�իVγv���r�N���S�Y��x�~�;@Z��*��GG����	�Q�i-�T��L��fZG�<�9�m�P4������
#�����&�.��_Y�>��-e��_�8�r�����@�����
��e`Ix�!����=�{Cܝg�ɡ4�Ư��j���*��_.2_`��k6�6-H��t�.O0���cLzRT���X�1	�x*L���E���쿇B�\WJ��8�0c����ùT1l�@�BX��C�'�w���9}���"��?WY����N��������g^��|���g_��x����5t`.'R}Ĳ�_'��[�=<�{��V�ug�&�x��ZI�A�b2F�T1���S��!` &?����%;�.��ԫH����y�ֿ�K0DJK&^����f�ϝX��p��1�͢wL�Y^TQp3������n�<M"��O]�,��@��I��gZ�D�E/�iy(�XO���qA�O��C!�u�F�7�P���������9/o)m�mC�r��׌f��V��k1=��ƙ�l\zJ���t$ f�[�-@3��9�)O���O@�t$h"'I�\�>/��н�娋)eAǆ�&��s���7�t�݂�S��~���2�HM��-@�½���ofy[��F���ˁ�M)�od�,�b�G�w�:֞���5���Q��ұ2:2��'�z�_FO|�LCg*���V�j^"t՚�z��b�\���Dn�o8>��O�����\���H�n>d4��a���m=+�*���JT7%�[h嘯��3ا&�(��G�ϐ����W���r��!�}f�J�.|���=	���	����M���������]>�����������H3(�-�Ĵyxjᓔ�?>B�j�Ki�pb�wx������#�)��qU�������<�;���R0D͵K(̪xQ�*�4�Y���f�l7y5x_�Cͬ�θ�*�lƗ�����o����lR����V~9+���e{*�|��,��#%9�?�Wθ��|.&R����5��%��%�_�����M�񁀝JAa��.(�\�= 4	����)APZ�5x��	�:��s@/����I�|��?�z��hl� ڭg���w�գ�� ;��?ƽ��g��O�	��{�ɘ�W6�ҭ�T~�t�˽d���c���w�0��d	@�񛐴����(�j	[�p�����'��b�;Y�Xz��S�R�Y���Ɇ�Ƈ�y�tp<s�#�vO�ز{�.6����{�\nv]�h)��?��t��Ff�>�UF1r՘TR>4��ӽ��2���s b�}*ֶ�y�v-��/�%��+r��ĺ�M7g9�-g
�.��l�$����Ic�&�2�)G���\Q�nq>��!_�8�>�� h�Sz��\���}�V9���p�{�+��͚���/�(pr�R2+�&z��NBh����doF2P�����)[t��Ǐ�Т�(2n��~?q�S�Л}�N�W4LU¬֩�M�(t�$��	ڱ7MH���t@�κ?w>�i)Պ�!�=�ȺA�� ���G|(J#�3f�kZ�|d	7�F����|P/�bN���m��6:ԜQ�5�C�Q|����
�.��4�=��z�W�)�%ϙb���g�??Pa�@��K[ϡ>�T�N���?�PY�l}>�A��Ya��	?�D���f��	����L)�ݝ�1qf|�]�J:����ǽ�Z�8A�Kҥ�p4��M^tM��Qeە��YuC���D@LDȯ�
�3���na}.��qX��^�{���e6F���Ѡ�n����Z �ұ���aNGe�,�l]�3�I*�L�tZ!EU�)��j�ږAm�\kof�yC��v0^���:���
8���'����r��P.?�`�z�5�2r��8�|�h�X�W`�O�L���N��/�Y�1G�c��8��5*Jж.�o2As F�r��|�vCY9��J]������oa'Y�ڗ�-��F���ؗ��{(��`r�\�AK �o��S4�������KE�\g���%ꨝ��#ފ�F�wIK��wo.�p��b���_gY����ˍ�����-� -��62m��E��k�?v�\�P�j_՞���u(�#��a�K���a�� ����8oUVz��T�t���ƭGD;A#q��0Nr~y����1��=��@X��*�|�U��+��y�'m���y&��Ym�����N�d������C9Z��j��aI����O�y�7i�i_<��3�����-��{�ﺍ�2u�jb3��Us<���c]RR; �H~�#� 7z�����-eI�ϰ"�?Z�޾�l�+��b�/���ђM ?���һ���V�ϛ�C{)_��E�l��F���}SS��!�do��zA��w���{{�:��|��գ�]���E4i����dkK�/�3��7��VjK����؃S�6E��{F��?v����{��YG��O��n?T��"'��2�:g1�g�	��.Ҏ���-����<��I��b^5f�g?;��e2	IF^�6x_GV�]��|��i�+�O�r(��L��[�$	yc�Ns,Yf��uh���$0:~�N����G�܏��J��mq��[�<u���Vw3�ր)H�]�����f�����%ej���h[Ȕ�O�6H��E��t�y�l�M��Pz����x >-޽�����f}T�-�3���_�����]	Po0����ħ^�fI�-`�����M�r.@YAY�8?����J�l��0^��a���3G��壔 z�N�,-)�WXԿBR�3��t�*S)������IyᴸD�`��dh�@�
��	�o|�y#E�g�kH�T.�	G �7��7`���0b�����~����σ2���k �ls�����kx��t��@�d�-_`F�p�.׆�0��>�+)\cjM��c��g>�V��V�ҶOV4�-p���Ȉ	q(�]K�e6��[rU�'#%�I��Ɲ]�֠�-Hi����Y�;;�֑���� ��v=J�Қ?�`����H�����_�[�� ^�f�dj�X~���*��˫-�}����׈�%w��x��`�-B腏h�?;�� L��r�e8);��T�3�)0��� �
�XJ������4G�ϮO��O��F�7*��#�v&�C֍�1G��KM�݁خ7i��(�0��('��A���Iј�rF�5F�&!)i*�`�Z��R9�Dl|�@,x���?�h#� p�B�Z�y	mR1�B]X�|?]���?�l|͋�5�S�|�*�(��/c]�!'2���b ^lpO�N�H�ԡ���G=�s��zL?X��;����e(au/8&�>X���d���I�z�Ĝ���ۗ�YYibD�4��j|j��~�����
�������ꬸ�\��,E)�l��(�^p!<��
Xc5\�f��Y��&X�H=s�M�̹�R@�3��#�>������?��!p��v�:C��*P�φ�4O�
�/�&��Y�X�Hp>���x�й��NH?�G�oC����ًk�B�U26/�DZ��o;��쌚��2���2���#�M������w+���66��r�ۋ���T�%T�p&H�XNR����u"��Y�[���1���o�8���*ٛ�o%y�Ҏ��f�����B]�wa�4!ّc�[-��\���xzHV�y3Z5nx�����k�R�v�����e�O�w�ha����5��a�܉u_�.G&�>ܕ(��+��F3ntym��� :��m�20(��M�s��\�7h��V>fw�0���HcsC��BhՈ�.��[�	Y���qa��"d?4�&T�͹�z�D'1�Ls��m�	y̳ܚ���Tz�d�g�6E�%ҏמ���g�����$H���f��vee"�� �����tր����KA��7S#y3��$���0��!�ɿ[>���d��S��D���&�W�K�>�m���ŻD�F �u�1�9Hy�'�V�$o~�yʵ�Ñ���/s~g�!/�>u�e�f�B۳]D�'�]�iM�����C��!�jݗ�^qӶ3�U�C�i�L�*�|��m�U�i |Q{�؈jF֐я�������Z��i�0����ʏ����jt�����4�3O%f<�Y����ݘa���Jc(�a������s�U.�tx0$��%0�����_����7�	����CM��T��t�y;VY��K��5E�5��=�6:�LD'�}���F�g8�Ho�9��Ğ��a-$r/���߯?��w7���9�G(=\��n�`z�G���=�S�q���2b����L��E"}�b!��:���-v���V�^c\P{$f[8���!��$x���U��Z�0� ���"+��m����KiQ	+�%x����DvX<�\�`��|{��0嬐R��ۡ��;x'����s)�ŹP�
 �M)/
<�a>H-��m����R�i�lH������p��Slv�+�c���k�8N�J6��Hd7+�v����!�>|m�J�:2���ǎ� �q��x�!��x�b}dD#���jVէ���	�d��hC����[KDf^���s�3�z{+m���H�j���%�a��12�ze���������)$���'F������٪��m�sY���j9,�R�J� A���㑴�E����yK;d�����Aז������1�w��gy'$�����������:;e���V��8d-[�1��Z>����Md�ac]:_|�ԕ���BC#q�tG��4����_������ɶ5r�\���1��N����O{�,]���b>���k��v���6�m�lT��H��{[�j�<����8*W�0�^@h�M5s���D�Jg���
�~�kP~|:.=iV�㛇��i��B!��$��m�<�Z1a}��#���iV�z�d俨]A~�X^���n*=JS�7h�69ؘ]T�i[�5���������&�
�i���B�b�#|~�5��|��!&���rM�m���Ws	�H�B�ꩪu�Q�p�]��Jbj�2�H<��#g\��=T,�l�
�!+����p�F��S��a" ��A�Z����0.�c��c�h�%��'��=%%t@����s�亦�w��4��iʩ �{���l��/F��݋w��h��+�!-"f].���tJSO�el� ���vM�
%J���Ϯ�S�vhU6��ת((e6�j?��}�[Y'� ��~.� �_�Kc�t���*$]��p����j�1ے����W�gu�R:7��9�^��B�����;�D���m��#���+3�$h��ߍN�N�D=��Vk5kܫi�%��4+?=�������w�|�_�AT�@����|}`��{3��槱q������0�2����_ҫu=��'��&�D1!�9�����
��p1~U����G0�[h�SU����D[�"6��-�3��$�{�Si>���y�5�<��Dh��r�Z�PaS�W/�h��֫D����E_<�$���Iۯ��%���o��-.���x3��j��Sa���R�qkxk=���{���#B؜�1h!��/��#��bD����LN�4��q;}{�4�ȗD�C��#�8�sc��w�Ub�0c~\10Cu�G�,늚a��6�+_�m��u��%���bzh�w���:.f��!Q$[�Ը�1�@�_6i1L�y>Vި](�c�Ւ@cH�Q�W4(&�[�'P��rss�v���a����ƫ��Kg���	|��%R0��.5��mՋ���Y�[���@6 ��xe���Ųe�h�p�q�jb'���؍|D�n~׎�:J��Fx��7n8���m�w�ٹ����=��h�U�;�J�>�$�JHQ<�Sئ�tT�g��
#d�\��6�ې�=����~eD�N�7���u�ҿ������"#Nh���E�ǰ�m�7�Q��r��?���4-��n���H$O�Eg_���"ѩ-y�>�<T��=�SVݳ���J̟��{;m1j�����'f�~������5����X�i�v2�X+�aVE�^�����&�����%.3��́�IL�m�U���ۿ
���O]��Y6)D�i�sr�i2r���rKJ�!uS���C�a�)(�AG ��oV�WVU�2*6��A+�މ���tɤ��a,gK��QU{��<jw�~�f�T�ܷɱL;pR)�W��4�QGo�g�7�3�����e�Iʼ�Mqt�����h4��K���/�h����.p}�f��H��q���4/�=�纟ݣ���~�ގ��+eM��M�A|<��9�Fu0+�#��$��5�t����Yso�M�XN?���5r���M��	�'����	��-X�웢d v�a�An��ӟsw��u����B)��(�2�s�Ҵ2Qo�́ @�]l��j�r��_��&�kvΒ؆�ǖ��ƣ���Tߒ���E'�&ٝK-X�O���.n�r}M�~�C�o���8���-U;��KKf4����ի����4����5Be��:k����8k@O/<X,޽�{}{��c��O�L�\&���v8W>f� ȁ��ш�a@s�Ӱ���Wt�lor����������"��'�(r����k\H��&&�İ��ِ ��Z
'`�^ĵ�H�$�U���O}��\Q\j���4���z��,[���	'�����u��%�	���וN/ŝNOy��7N��e
I�&#t|1����S��`|�Å?��Bhňt� �ᡣ��6qIt@f!�����^���0�����H�2�P�r� �d���HD5��;Ⱦ
	TEQs��$��r�'�n$ޙl3��u7�FūQ�����T���܂�&{7T��&؆j�N��
c��	j��6.��
��r�9WY}�C�<mK���8T�n��J�(��lMl�T��-�]���vC�����U�r:y+��a�xm�BBf����ߡj�HV&YD�~.
�w�������wB-�����ؒ<_���C[{`m����Uc����n�X��a�;��
�W��A���V^�#l�������>.�C�Y�I�/��x�a��Zʷ4=v8�FO��A�GY�1��J����R��dZZّyS�,1(��BF@l����P�*� ^V������R��G9gLOh�'��V�o�����Eup������)P�IL�钌��w�>O3+���]�e>�^m�N�wƬ��*��B rtY��J�E4e��k)R�Ζ� !�UƵ�f�B���^˳��B'����_ʕ ��*3}��&t�~-L������Ke�`Qҋ(M>X,I�)
)����P�}�\�q�zL&��u�q��(Ж�Q����qq۬����-E���z	|t�yq?C���a�i�Q:��C2��b�/����沭*��'l >50�-�f�=_�ӳk�s\��q8�b��o�~*(�_��yI�M7r|��G!9��k�l�����RR��Z~V د�w���x��}��`����FX�G|�� �k��ڨ��̕u�	����J�K� �J
f�p��#Q�quX�T�T0��︤e��pd�6ϖ*�	MS�P�}7٤�rL?�B�[[��\a�scP@/ȋǖ��zo�Ƃ�q5c���B1+7C�ls�Jnĺ�q���u�<I���Q�T�^���l���SF��	���UW�"��TC�t�����#��.��T��z#N��,�@j���d�ɑ?̓h٬cv&&��όai��o�g�+A�B=��԰=�Q�w�ǧ�����;p��M}�9�4�87�u����9a�,���㠃4v'�0ӝ��|kEѼ��2�"g{�_9�����'�[���7���	c�dS�	6����W��ܔ,�\q��Ќ&�i�2�&Q�֚���@y�M�0�Ђ+}.%xM�U�<�2�����'�l�,JG�M%V�|`Z/���-�9r뉺���Q��oc7��JJ�6 oU�|(
ю,��\��	8Qah�����t�>w�� W��0���i������V�AڰVBJ��T���6zވ��ٖx�Fr'�행�y�2��:qbh7ʖq���n�,['���S�𔉶��~����:�E���tM��R��; �/��j������3���ԟ��!��
�,���z�q�t�R��d��Qj��f#Qz��}껐��B�lװ��~���ۉ7���l��u���W�N�H�V��-��R�4T��ʛ5߈��4���
�BlT%�sAtgZf�E\�H�~��V���_/Ճ��6L�:7c�-��W�����L�
�c�>H O'%e0���*x�d0�%�Bs*���XMC��_����S�!%�W���{4�$X' ���R%
m��S�����(Wޝ6n��`eO�E��W��.G��3*�3���mC\���D�L�%�C��l�;�S����MBK%Ѵ���(��4�S;�QLk����J
ĭ:Ԭ`�#g���jUfv���%:���7B}A��-���z)oLI 3;�$���_�~t ' �j4�oMy�V_��Y�y�Y��C%\L�-��R�3����sx5�������H�H�T�4\��k)��&�x���]8�,�����o�U,����* �u+-�?�f(cU�R)LĴOI��L�!��u#7]]u-o�9=��M�+;�)�K���cQ���)����_�]A���ETi��?}rU2J ŲE䆸'�L��ueM�_v��?�}>�H�S�НX�0GM�6�ureQi@�� z��;��ǣ�.���V�͛��D�E���9%F��ܭ��|��6ڍ���be<�$$�_�+��%}�gh�I@�9W�=�L�`1sS�X�F�%��.�����Ա�?)��k�~�u�Q�#'?|�����Ey������`��1���k5��O�d2�	6���[��O<d�W� ,�!��Mx�"y�oMF��u��ƃ	jLX�b�o/�P(;�B?�u �wS^5�O3�f���E�h�_�.>DX�3�c�
ȤIP��n8��Ƣ��i��vc9ʘG��%�����)�r
���$Z��C�00}b�F
�L$d �M�#�kl���3����0���O!�I�ɿ���j>T0�%�fC{^mM���b��h�3��t��Q��Ŏ|֐�oH{z������W��x��"����f2�x�i�h݇Nܳ��N00��3�7��P�@y���O��[��tT�,����yP�?��i��%��W��:6��H��:c�?I�2�����d�N�Z ���2n��>m�����j#���8�z:���<���p-ϯ�a�Da0�)N���������ҹJ��d����Gfw�T��ߡ%B�Y��GI��7����h����=j�R1���`6��6�*R�4��V�,���!�&N_�c�����N����Ǳ��zNK��.��J1L�k�	ȶ�B�t���*qnb`�s��>�/(��Br�Ԗ�.QǔKmJM*�`�<�ѥ|��,�$�V&���?�Y�̦��b߻�X���v6��\�30�h�Q��vC|�<0���T� j��fP�s�m�o�D��h6�;G��d)�7.�y+�~�Ff=Ùm:Js�*\wٰ�𹹦��`Au�S�_yqo>�jXZj�~�c�aLṠ����f��|-R�A�
U<��tJ?���p��P�6��
kP��W
�0�%��"���ST�'`��f�l�~�V�~�X�<�Y��g�TŅ�ݓB�N~@#�Y6��&x�E򄔩��R�k��5kQ���_M(��C-��x0�J��Ӑ���}Q����6�;	Yy�~^�dkƩ��<���^����P��;��`w�� �qt�����h�:�e�*r��]��XK�q/�D^ �b�-�MB��/�5n�v�����*h�vp�&�}g{��;;3��:D�cCb(M�vBw�A����mõG�w�ЎN�oh����,��dl&�|����7.��b��0���`^������少WT	c��[ ���H!x���)/�]��f]w7�.O`,�Sj[�H�?ej���n�i�ny�SdKpȠp[Kp9�b�,¡�a����M�A�x��W18�^o)�W#ۤC�w�Np�r�%�:YX���0?���±��_;��0��ӄ�D���_rI&u�Q��Ⱦ"7�+�s���z�R?~�%O~剸��?�g�G@+mzO^B�"�ET[c�[6yZ/Ԃ�Oe��w�����Am�6�G@��6&�g��w�{�|ꣶ_�d�G���fd��Ȟ@�aW��?���C� x&� ,��Xs���O�,�����)oCM���Bj?ء�N[oMN7�J�F��!�@�8)�F�ښ�&�Y����1���e��^'�9�r����'7�y�Z��(�'8N�����졁��VQ�S4r>�2�=��$㎥�9���(`�=�~�p�a��E��2�(G�8e�"Ďӛ���'���A�"N{�\Ûzg`�dok�J�.�9!�Ojle������6�l�Ra�O�j� J�L�/=1ק��G���<�_'?�: �O���paS /�\��C	+?����{�4�Ψ��@��\�+���=4��ek�QJ;���z 5�]\&μ����M2N� C���U{�*^��
����ƢJ��@�C]�ců2�K��+@9����$��z������U��~P�w߃���� 
��8������j30Ji/�$���O�.��3�7�t9K��yLB���>u�w�x��}��Y'������^�)-n��zD�hh�qoP����Q&���
�����j��6��}7�o^�Pu$� ��4�p$(;nk$��y�g�e5�_P1F��?���Yx�BQ�����x�|�h��i7ω@H��e#s{��,;!*��2p���ۈٶ�������F/+J������W�o�:_q�����|]}����<<��E���Q�
�K��������.��>兡�E�f �$cw[� �Ñ�b���M9����dX�>e}��>f�� �4CWQ�yy$eL����[AAw<X`x��ƍ���#4 Qs��n���<�A]��]�QbB]��eP���UB����2��#tҡv�,D:,���@� ����b���$͑]��V>��#��WE�3�r?	�衧�v7Vf�d�#����f��z��a�bn�1�m�.W5�ڰ��'WO��H�J%�۽���?YiE����#��Jp����w��Nw�4K(���]��L��P���)��cٶ��2�ሩٷ�V�p����`q�1���H6Q3~6fp�����*�,ߝ���*��J?����}�{�����������:���-4�`�GA%��C�l`� ]�]�e�����u���bS{���D@+ﻝ��p�-�B���n��<~�� �,�j�bB!M���yni1`�n�e��VOٕ-h[m^���d�O�B���ol�I-?�� ��% �~�6�9F�>2:?8a���\[�]��\(_B�D��G?�q,���	�ŦcW�-q?
A�ٱ��D�a���I�/ ��m�fo	`��[]`i���+_Y{���� `�2����V4�l�T�ذ�j��H`+~�ܳ�U��*�q���ss���� #���]�_��n�Z�� ��9/� D����l<S
���Ɍ�M٨�	��������փn� �p"�8����@��<��ĸZG�w��m��"\]�3��ԁ�w�I����m��v٤�Ox"�*���yW�'�J/��C�]�A[��]�_P�R�jٞ�&��F���X�xֆA�ɒ�����[�@��Z/U
B����8d�d���G=�Y�LN7UJt@����
�fß���|�����9����2�J����%+��M����!�ၽT��Z�q������B��-�Ђ�����x�o����ˆ�����,���;FנP�g��cJM��eu���� ���{�xֶ39�FPՌ��Y���q����yv���nωH&�!� �w�x���樘V���4,m�\��Qխ�ɰ`/��<��Ǿ� �[T��B[1���BM���Ui;��mE2�]Z$��E���DV
>�Ϥu��8A?F�����ڟV���?����	M� ������H���Y��&��,
Ҍ�}8� FI������râU.�+�A~{p����r�7(�D�5۹��ԃ"�n]���i��N�]D�lq�ʤr��P�EǲŰ���坼:�Je��g�7Q�0V�9.-b�Wl�͜�ج:kѨ"��%��e7��9��g 1R �_���".M�|l��_���1""&���\1�WY���ڨ��H?��TΞҊ܋.�!ꮷ�ƺ���W9x>n��q��J�� U�f��?���v�2?i�K,1�=�A���O����Ph�F���H~T ��.bɂ���t���JO6�b]�Ya��+�g`�4�H�][��x�\�%WV�;��	^�m���z�ô����B�]'����wL�7���_���=UQ�ӄA�0ף~��h���k�+R_�,f�)�FCY+K��'�S�������	��R��S��&n�b����Q�Oꁕ/Ѵ�s7�܀�?���� ��0	�F�nv:���O#�j��t�L��a
�vSf�|d����[�,���>j�FIǥ�$����:��sDg�s�&hg��m�C��4o��m��u|�KG|��� K�BD(75#^�. ����&�x�ڱ�)��MưaTi���HVD�n�bXM#P�NA��DY����ahr0N��ʃ�a�R3��J��08>�ړG�Ҹ-L��(&���T֧��r��=��P�tWc_�E '��C�������3�XL�&���y���XJ��R�<K�j��������,����$��aB2:�	��q)�|a�#A`A��ɚ�4�ؤ})M&���L�����=Ѐjez�47BC+�I��y�3k�Ӽ�-�ve�h���?��+�������x)�B���8ln�6D���t�P�z:��sf�_/�}u"���?v����i�P�ޛmҌg�/v=�O���ooV�ٌQ��D��h��엮�c!�ڽ�Y���R���Jݐ��c���P_b���������㻔R���Iá\�ŏ���?�"A�bG��sTo�CW_�}Pp)<�?3 rC���([�8wF�LQ�	M"��e:�W�
1	n�:�隣t�����@�אeh��Kc�������$	  픔֟G����
�ɻ�
�ꏕ��N�IS�U>R�5+�\-M�'PIN*��,���HZI�U���eg��新|����K.����D�D=����q0:�)f\�RhH�7{_/�-z����ƭ�*��<7t^ί]�U+��3�B��C��EVe����6q<U,��Ȗ�KU�U��|j�׫:{����J���@�
� l�q4b�ڳ��X��%�`q8��7�|�����#R����4*!&tD�?�	����*>z{�#T��ҴmC�G`�>7��P���� ���!Q=��y�ۜ��'*���'L�ɓ�6�vq�$�5o%pM"�ܛn�Ŀ�����S �R��@7��[�����|�,j٩��	)�����n�:0��@�N%�G��6��hP�$[�q3�O=��Ԝ�#]���\��t�*[b�t9�L��p�*�}ڿ�"������K�s��eDxZ�s�VҐ��<�����?���DX�)���	�[�Ýf�'<�,Z��lb�L���� �#�vj�m���t���{Y�sf��XD����l�r�w%��4��N�?#5���r,a���W�YD�e
NIN6���D��V�@WV���o�5g$���	PK�eo�Ђ.%�V:̲{Q�KԚjr݇F|��	�_~�NKʹ`Ol~��{:�[�x��Vu�J*S��<��:�-������9)�jF���Pj��._���u�T�D�#d�����/�f�ȏ)p퐗�+P���p���}�?r֞�����i�<��k%a��p��G_�_5���~c6�R�iFрL.����r��dm��ӊF���-8��xy

3G":W*����i�0?g�븷sEns��A6x�}v�E�
bU�4?)-c�ல�����8��`��7t�E�U�'��,�����*�̷+_4����#ZZ�s�T���J84)���eOb�~�%�#� k�U�Y�e\."F��}OR_I��Է5G��S��(�6��b�\{��;���Q��t,+_�}W�x���,����<9|L�����ֲ$�+�B�}(�Er��ϡ	R��]�]����g,v�ܼ���_o��#�,�m�?�����~b?�7�����~�|�Fc!��asm~�X3��H������	J4��°GH��L�Op8�
��n2����0��9ɓ����ݐ#���B���^���+�eІ���9�"d�Q��1@y���0cSq���<]^"��c9Fr�M���q���c�u� B�bd���r�X��-*�(I�
9"?2���:��>�K��#W~�C��\o��/z�J���R� ��1���4�X>H1�]o������X�u���AԽ��TW�0��L���j��6����~6LTC+	��K7���A� �p��WC�q<К|� 1�H9)����e�	%��^�ft��RuH���$�^ʋ��-�
Y�Գ���4R��[!�T���W������:/#��?��x��*�`��7���4��s�?�� ~�Uqo{ښ���.�'k�r���9ז-��M@~=*'�幢PH�O�h]�us0���G,�O,�t^�R!�/��[0,QC/R���F!����b�:` #�E�뵤N��>H:����b�9����v�d��}���Ӟجy�q*��$Ps�n�ǠZ��d��{0½_�r��@S�lGRۢ�&�`�
�U!I�����6jK
��݈��B��<�f_Dڟ�Gʋ� Հ���u�7)�y�#Ӫ5���ДQ^	��b�T��Ym��fk�N�����f������J�J�-�ހ��*
�߯i:��t��=�1�j�]��&pH.�)�W� �ۯS&$��C���J$?ԗ�op(�&��P��ۀLz���?]����!��]zi*����ӥ'?��W[(��������b%!�.���Wt����]�)�����n44Vٯ�v��{��@=J?t8 D	�*�|�|Z�}�a�[E��MO :2�8P'���ȕ��ҟ�<�y5�Z!J�߉�Z��2K���s�B?�;;��sr#���A4�)�y�1jO�k���k��n,50�]�ߐ��c����0�l�j|�Zc�	���J[�Z�j%�p���#��|FIy�Z$a��&��[e�j��ݣ��"���j1:�Ss�SU�:�g�D��J�Ҹ)R��L�Y7Vtx�|n�k�P�;�#���ؔ��Y'��Mi_�i�CH(�f�xŅ9�����ST���g6UMn��e;��vC�;b�	ӟ�'��`��Hq��z콣����~ �+�u.���06d�)��C	���.�Pjnx�.89�:8k3W�Y�-)o�zL�%��Wh\뺰��Y1�@�Z!��q�
��8tI�����_�V�D`'�]-A;�0>ǽC�~���D��B�r��[x\:_F��1q(G#{� Ҍ�zp�B��GG�O���ϴE.pQ4��QQ�D�7F��6r �a�o�96����X��&<�Q��L�n[�kդ�����f7�u'Qk�@�3w�b�>(��jp������1�ҧ4ʫ�C�����c�l��-ـ���f�d���3���i����9�)�Te�g�0]�B�ү2����qA�
ꛦ|�#�V�/O55�U7�"�G�'E���hsÏ5�x!�� ������8\O��@���I���6�</�-W���-N�{?�=b|6B��RY|a�N��ܖ���l�`?�`:	S
f��g�>�s� A*f�ǁ��s��P���~���M��DT:�vX=RW�P��%���׉��,��SnC�qÙaL�S?�̄�d��7����g�Ѵc���,u=�ϡ�ZEm�&�����3�,!BW�*Bw���S���|A�iC5��h���͘5�r�WR^݁�}e�Y��*E[$+Ou�ES��aUV���IU>	m�LS�J�w�׫����`�{s^򚟴RA�Hb�DsO����oi���n���BY0i���?)9�a�8�/fV$���8�:I��ЮZ�d��	��퇨��U-��vR��%�Q�~G��`�.]�L��l��֩a�^@-���K�������I�BR@�sC�t�#��V�@֕��`�J��|k�d�ݚ$J���K̯{���.̠�z?hgA���"e�a��o h�.�d��u5e���s�!���K��}̝I���g�]_	.���?�"+L6y�Y����lN��v�9�� @J�_qcF�V_���S��/&8�K�i����.-��B��Y�����:�� E�G�`�N6!Bƣ������;�>_��|�c� wx�VI� }�M1T��i���ª[*�2�+�Ϛn���w�dF��e�%'��?�~�Z<��P>gр|:ya�5�Zo���Yld����K�X����/Pנ���AojG�C����G��I�^d���o�ԍ���^�ZQ�q=��)��tV��[�^���}�����0j 2��&����k���Cg�Y�0����<)$��l�s�n0vz^�O�*4�\�s�u���>��:6�{|퐫pŜ�qU�ls�|��>�M���~�>E��2��H�
0���C��!h�?ׂ�4�`��0�x�9�D��a�"�PJ�g6�U]��_�s�ߺ�����^�vB-����zFz.�sd.
�F/�������b�Vt
���rS���(G.�!1sշD�:F��n��bֺy�A<�ǰ��&K�_�.sG�xz�1t�E�A��ŀ�I���+�&���&`+2Լ������4J�[m�ۿ����4���\,�ܝDm��n��䈈z#�@����K��`XS���s�Skp���aW�.~>������=�D�B��YmV@
Y���<#�:��~�w��3
�|�vOH����D�����l^�g?���t��kL������m�S{Ν���p�\��x����1��}f�"=��3Qۂ�z`*ؑ�����(��R����	�qj��Ԑ������j���;��w�Na55� �tX���Ћ�{���ڍd6}�"9=1��~��S�%ain28��ӂ���	���`�|�Tr�S��]��?p��<��}g���-���7aw�h0�S3${R���oo���~8EB�� *���EVv&���ق/.�*s�sg�������!^�*Ti�zK+�C �Q;?�dĶ�Cf�ˊ4ݔ��J��w���^<��]"Xk����u$]ںM��S��CB��&��'"vUK���C�@�C� �qp|�!o��2�2��+�3�9a.9�a�J��]�:�E�]dӊ�h����5��`i�������eSj<�@��Js�d�����zRž6!�?�.����!��< �qj���h#\FK o�)M�����`Y92�{�I���Ob�$�h��z��Kn��.�ڼ
��?]8s�E�����;�CL�����Fk#	&��}3����;�)�/��4|d���g����39nHY^D��C]���l6@�/��U��yx�a�/Rj�Eo@���?}��
 7�Ҽ,w�x�6�ص�4:��A���E0Aff����-���>Cg]��\�b{z&e�T��5�|K/����h����42G�qrXja]�"��,��1�:�R�����SuJ�ME�c5�ޕ���t�If�������}ߖ�������9E����y�+�H*~���������X�S��P�8���j}���i��~����/V8X���Ơ�u�"k���+D�i�����i8��Ä]
j�z:��tb[@�v�R#S��CIn�����N 2����-��vu�Sِ|��y�����u.w��p����K&P���-��"+��W�<[[�H�	�	�r��lj{���g�W�ka���qw%:������
�qy�,��!���IGd���[T�}��o��
���k�2�_e)F֖�$ı�=�w�ߜHʆ1����@5����9f���o=raK{�r�ow?z�{D�.�o ��5Z�,�fr�蓺2|�[���l����O�S󚒍���Y �ą&�r�_Q_��U������H��b�p��_uyxB��&$�[�ao�	�c�"��6� I��S�3�7W	��K�
�*�"u_>��+?��-B]��{ܑ��n�B����b�Ň��+5��K,*<�+-/V(:Ri���|����`�';|
K������\���?���v�6��)�Ȝ,]�A�M�8���G�<{��$�l)�8�k"��m�^���G��Bo}1*X37#j�Q1:��-ӈŀ�?�fedY���bP�	��f��� lgڕ�~�����*�Uw40�Қ��u�gzٗ㠅�H������lp�sɵ1��e�/��CQ��5�/��8C(m�Uݞ��o�מmL�F�*�c�Hm>�3���ˡm0�Y�w�x�`�'��.�=�#�߄�}-�IA�Q0i9�K���8���}sETi.��i�y`0a�|g� �9��љ��i#�]3aZ y4�8�'��؎yYm�$	A:�zv<���	p�EH\��#5��GL;��X��㩕��o��T\��ZB�)s�ʦ��݈H�� U����W�ᨮ��jr/�t���:e��ђ�f&���V|��o�#����^P�\�$����^Y �/X�L�o)�X��O}ۓ���X��8�U>��}��MD�_~������-3�)��U�n)���k!(,�B������8�2*�X�!ܼ�j��Ɩ�j�Ԫ��dh<W����?�d�c�H�=��Ꞅ�Y�������h�݀�L���I2�eK4qEm��D�3ض̬B/as��/�vh�d�)�`�:� x7p��L���i ����-���{�\ה{PA���B�`�0���0�ۅvv\�U%?����yϾ�ܳ��C	 D��q�K����ucX�1�\���vX
bթ�a`��-�噤3h�Mr�<���8S]}Ƕ}��+8���.�5�����ǥ���D���lч�D�4����U�!���H��_U�V/�*0:�pZ�[#
Q���>�Ĵ-�y�	\�]歾�=W����=�*'�Z�y���w[ĩb!l�;���y�R>� Z�R��W'����Z@�SG�f��E�����:�Gg���:Rg���~XSl>މ���tw��Sn��ݘ�@yÆ�V�N���Y��g�W���=�$?
�i��W4QEkM����_��T�V��H(qvr&+̚����f����E��t�"u���G";\
S���n�ޅ��x҈h���y�ob���Y�������b��u
^e����SoO�b�_a�^�˹v8�9��x�5 ��K����@	��3;�zP�.�|�����Ȉ�r��Ï�X��tA����d�R�Ӊ�A#^	�Q��L���|Ʈ�o��� &�o��=�T�4���8�Sio��9N�r�&(��`�ȸ +2���0U��R^����Q��za�RNG�k摿ܜȆ���;;o�o.�K���D̶�:�/w!����g�����#��U� �!R�ϢT�M9e>�e~�@�"��`�8+y�,gN��n{�q�G�Wԫ��:��ф��mBk8��u.���ĂI�8ky�R{�ǅ���k��Čq�4���1��d^OIE4���b?\O)C��G��a���F��� ����&ER�{�;�����ÆL=7�}��s-R�]e���iSF!T
�Ҩ[�,�X�
is�X9��?c`���#H��F�ߙ �2|X��|��Z�����2ӌzF吘�
��LmysLX�,qrm�Tk�w�h�Ӥ��s[�QL���	�q�D��9b�
I`{�l�� ���,z�(��/h�1E���+��W�쉉�/˫��}j� p��y ���9��\�؝=��Ջ��SIN
����$t���1�u^��GÅ��X3�}�Q�\�w�bci�( 9��CNg�����ka~
L-�W��[n���,$�%H"���t�RQ*܎�����v��="֬MJY�����9i��f`���]�<s�H��"Ec��q�;������ά��it�v�[$3
֢c3��m��i�*�@�GpbBR�du˫�J_Qt��fՙ���'�_��N����p��@.�dT�G�c�F���u8ĸz�%�ê��y ��d�vhD��U��d�����J���R?ȟ�3�#zi��]���H)n(��C�aX�R���*b't*��[���J��a�A�4#�}��e�_���M����T>�ݝ�jv�t����l3��@����3��ɢA�z�D��H�+���I���n���ԵraFٳ��$�X����I�Q$ZQ���Kxmv�'�	sW�y�V�_-�V�<�mHֲi��rs:�L��8�[$V�-��R<�\޵As� �[[�(I�N�~� >5�V��ng�?!�	g^�{.>�qh�'��E���y\ĨTߐ<W(�� ]Z���bL<ur�#jr*o/	�#�9hvs���&��J(Լ�Fch���)z��' �Ws�n$p;\>(�.e�e�*
9���fԪ�BK��q%A�NT �Z�+��±Չh/����n횃����&��V�ڴO���`�VWM����5� ܝ3Xo']в\÷��:�����х���[b&�nteG��zG�91)��Z����xӌ����qk=���"��Zb�}qC5Vw��4K.^�={��U��@4�x5�H���V�X�3�65kԋcmFRZ���@-{��rGt�CQ�kFw林�����;u'ߨ�c_z) ׬�������z	;S��xc'�Ϗ����oL?���m�|���@��0-���LS#�M�NW8��*�%.���կ�Q.��R߂�הqnяD ���p��xc*c�U��l]����.F����O��X=>����1��#,�O@��pߔ8��$�)4.��ц����;��'��*2~�˚H�ȱ�r�f� L
��(ty��q9�J Ax0*�����mC�1�V��z����1�/axR�� 䩎�#�CP�F���ЌBV����k�FN,(KVJmzl����i������Sb�g<�{�L�������_� 1$ãvcd�ܕ�������/�V^a������;a����Kq�u�5} ��Ќ�>OQ<��q��0��ӇgKL�nP�3����:A\E���9��f�U+�DĄ�due�}/m$���x�3�
O�s��4�t�W�qLm�~�2�o@Gl���3���������cD(9��P#>��u2�j���X�-H��ݢ%�0��ЎJu�%�H�;l���X���%6yŧK]@ ��P�{���K�#λ T�Z�������b�ƹ����k�*WfG6�=Qu8�KJ��yWk��gxl�l0ԓ��y�w�bc~�Ӛ��;�Bw�`�0P6h��D>W�.��)M%B��dG?��w��Ɲ;d׋q���V��u(�;U*�{y`\}jq�c�TҠ�����c�NP��W���`��k��J.�Y�m�ͦ��� A�D�a(������GM^%�,��X�:e<��|�a+vtjf������(�I~����UdN��tfA1�[���9̔n]�oQ�H���"Ț�?~�0�K��ח3E � �mq�K��A�� 0�;�p�U�^B����s[�Ȯ�4dY/� iX���@dN%]�[!�9%`~[�2��H��t����=���Y{-��b�R�-y���H�����w0C�@�l��Q�����n��� t���ȶI�v��r���M�aKm��Z�����篏�$�Q��Q4�=����`���e1�u�$�#�ω����TWF���we���RWX�>/y���I,���˧�ZU=�b�s�������[>�=�ϼ�����(�w��ON��I2_�����#4�7�^،��V7��miÃ�\Q��:9?�ʗ���A�����;�s�.X��صZ����1Ҕ�8 �g�F�F{@ "#ɷ��ԏ�����%�c<\t��AE�N߄ZJ�^����+t��z��V�B��ۥ6�����A��@&?�����K��R�D�D�3��H9ۖn��TZ����f�=��Y)*}�>Y��R�9������r?R%��CA�A�m�K��ߩkP��q6�Z�A�*Bk��k���T�g}>��@|=$�OdN���R�!�Q��-���]��釛E�|z	;'ؘ$|�\j���
1whk֑��a���|���z(�ӌ�dտ��Z{��K�f�O������l� 1��.�(�	H��Z_qvcy��a��tĸ����+��On�� _�q�Qa�8�Ʉ�sE�j�k( 	��������"ӆ9Kft����p)X����� XLK�ɛp0ƽc�T��Cv�2#.������-_����\�W�ܛ���� �&,��nL9����n�ܚ����(��P�2�N솉E���#:���}`�9�ot���q�K�=KK\��=e��8LkX���~ʻ�d+#6�-ҿ"�5���,��OK���f��^�`�ڶD�C�3�r�����\*`�,,]K[ކ���ؙ��	�ş�<�6SXۜ�#�8�\K��������v ��詬��H��	e���0��+��DG̙����qBq��)nY:Cd�KH�����$Û�b{[�����+7�q�I�A��I�-��f9��2��,�q?q�u�i} �vmpZRp5L�p`I����>��<�f��9NU�w�OW&�����0F_��Ҥ	u�X�3�ZL�}E��ch�R�%1֗�g`w��,��h�����XqZw�l:���k���ڴI@��E�S����?+�>��%̿5T�܌�E�Z���tm	��U�w7G��� �41��4ux�,���`�Z�`�ͷ��*D�M}�"�X���ߍ8�G$��i��V=[�8�ZC��@�R3ࡣ�����?׶�qD��}_����A_�'�3�Qbq.�8���k�o�^��|̃.k���O��|x+�}�w��@n�)g'�(?�LH�%7j�9�GlK�v���ӑ�H��]�ucF�a���S�9Q�U��%��S�Z��v����U��ͦ�K�m
��~�IS���:�Jk�r���=�a�H;�N�f0z���w7O�X2�u��vц"�fkX�\KR���g��:l��Ŀ�5����e9�1P��Ve�KU�����N�G�q\=����{"J�ˊ�w$jgh$C�fy�8�lS<��5�aGOC�Kz��I�%v�3=[bhn^�r�'
юkI�u+K��g��LB30b4�ŏ𙈤l�S��4��6Wc�ۡ�4
���[���t��G2Z�	�&|\��������0w�J��*��iF� �P��2��k���B�P@���O�̃}���e�ؘ�3?���=�,0�����:�����0�L�]u |�#�+.�sS�@��%P�eRWG��wHO��Q ?������ ��tPDO��1��2�ҙ����%�"�ֳ��������,C���\/T��!gv��GL�����-��i���2�:.r��A'���X^�*exJo�DZE/��+�m�4��1L�,X�:��M��ǌL��Tf+�e�Zb��+0�oWG20;�*?��D2����.��5�����L%�ai;W����J�٥�������֞��q���]h)0񗤗�=,i�fu�=�� i3���:���24FQ�]3\y�gM�g��jF��Q��X�����H19\�u������\��㯓:�o�|,
�/o�-�~[�ؗ!���D��{�?{Y{���1�i/���R�^�қ}�0���`����\b��=ΉS�d�����sl�ַ��/�9���a����#ɞ�M��+m�΃��X:.@�����bs���=B��?Z����1��v2��/*u�\
��Y�[Ok[�����hl�*	���k@�DǤ�@��@9rP�V��'��-����~�M߱u���2�'�DS�<�ND<�(��Փ�arW� �<nѲ�E�J�#	��r]�HtGz�)�ώ��wP.|y�~MG���-�?v��[����4(7� ��lmz"���7-�m�T�pTSO��(OD�yp5��ӕZm4�x*��^B��3+|fø)u���'2���GpD��Sx},��E%Vs�.}!�n�X��9�e�)��@�d㿡�z��rc��A��<�K=[8X�MÏq.�,H+��O���b��,��D�jIJ���eة�Y1�I�ۼ{�Sܟ����W���P�f<J���	���9:�#b�p!|�$T8q�WG��L���>j�w��m.��0��u�_��9�F+^����hX�M}�o���~6aQ�v���(Si�\��hN����ê��p��z�o}�ti�����5H���"?�('���]L��?���r�m���>�R�`��>_E�Z�����!� �2���l�Hk��r�}4�p(���p��¸�QT)�*;Shu�i�,en��A_�u�����L	y܅�(��"+�
V~���{����u�V���>%�X��*���p���X��S�BZ�	���"�F�E�Q�1oYY��'lJ�����
P�jj1(�����. G���<��AKYY���^E���t��s�x�{Ϡ�-�e�,��i�׽���>H��D�2v���jf��2b�3��}T����06*]2{�iӡ�BD�h��el0�N��<� #�9*z�Z�AC��2�dѓ`�����TU��-B�̈�y�w��^]�uڵRk)�V�˅��uk�ފk��w�n�F��X<,�e�����9֩�7���""����:�^>�#�UN�a�����v��s����7Ԣ�;6�w}�
 N����z�c�[���(�x����&��fk&�'�?��$9�9�Wff��Y��GCZ�;Hv�f�I�l�*!����7h�|VC�0����W��+E�^C�U>���z�K������� u�d�F/$	����j��P��R�W�Z57��^������-�g`�A^��Ff���a����k��޹�F��e���2NV�~	�@����:L�X��]|c8;����h[�XZw�j���`9���f3�\>Є��Op�pƈy��>�[�ڞ|c����קH^��'�=����Χ~�UI1��!�M�PT<�4�4�:��Nm�T��.���C�2�c��ܨ~��3��e�
e2��7�	"��h�Mx�dlJ���Ǻ��G#B��)_]�3�h�ߒ�Í5���p�b�TNR^Y�N5j.�H�Zl��S1�!.L�(����`�N/&D{���_+�$Wnd����T�9N�f��7�]l�bV�Q.��M�K�&�<�\)�>���#V��C	e86 ��Q��!mZ
��B�f���9�/��2N�{l�k�|P���t6��|�\��߰$�]�s�� L^�`�Rg[=@�ϕh�'�8s��>p[HJ0ls���:
sKN�rGZ�Q��}����ײu��p+(S �"�9��H��k]Tw��\G�*M�FR,v'��~u�|I��h��jHHU�jLr�+Ã��tp�+^�7ie<�Oi.[����D-�^�[�F ���_��
l��S�b���OXA�Nn+�}X$���o���upZ��]/��z�;	6ֹ"T	��B�N�;D#r����r�Ç����a�z�8gJ����l�̦Z���.�7-:��-��	�L�dn���s�7���ɡa5�J��hj�41Uc����� 0WHϥ�μ �&G"e��H(���ڸ�v�:�Yя��9�l�멑"#S�㦡`y��T��@�\!��f�9��_Q���?2�F,������t����1O9�j�c��$5�F�ц���z���f�]Y����Mx���-m�^��][���>��k# �F*B���o[eJ������Vm��G�~��\vZ#�ˍ7�W(o�d�-�+dR�Q9�:[�B�,"|r�����c�2���.����Ld5��^I��Np!��J�VU���)����H��u`tC4��IW��+@��s��5�Ɩ2Ug��P��3t�����<
ӌ��S!/�pVx��h��5ݟVε��
ө�4]���"�g`�pR54|ӝ���;��'#""x~ƺ%	>C!]�X�m���M����ː����`���}�������[�\u��|��@�t/�9�/��+}�6�e�3��ށ�攵�`y3Ժ�R��������pcʉ:�l�������ib�=���fb*��q�2��ⓥ�654�'P�lx�PR6{#�+��|�6OTr���ٔb���.�MOf��Ⲓ,]�M�u����)�5��Z�Us���>�6x�`�[�)W]8��Lz1�\E�}-Ʒ�8l���-��lB>��dZ�L�<N{A��՜��TNU�����B�ő��uD3�|�ѓ��9�G-6�� |#9J��Z����1
DTݭ��UQ�a5������<���h}U��u��K��)csEZk�����7j\�7.��
�h�47X0��7�@�ʖ n�.��А�i}����l�$���;����?�T���&{ɹN��	��P���" �6C���G��Р?��`�:~���e;������w��Z$X��#�کK�(Z��3++ŀZ�.|M�5��N���N��4H+��a��H��ûP|�ze�����$�r�<?��\�o���8J��A^h'����b��zϖ���Eu V�Jz�e��چ�澚4t y��X�P7?�d`N��1��{?^��頬�ٹ�������u4e�����з��"�Q�0�� 1�!�[So��O�S�k@���tc�q	��{@GRA�g	E�_ӯ&�i�M�u'�diw�����)�6��jS��UQ������z��V+86�׬M�t����T�8L*O)��}��<�	����DT98eRS��aN��쩅����أ���=�5_��}��LQM]����n&]a\�Z�[�x[��\��uf����N���y����Y,W��T�Fa�i@ūT��mK��Ev�a�>��BZ!�wF�[��+���m�� c��|�U�P�����^"Q����_ۙ����ش@&ҳU��deb
��8ย(����x��j�٬x�Mѳ�oxo=J*Lne� ��۞&Қ~�VC�P�݊GM���W5�vBWSmB#�U��z�C���.4���#Q[�fs����a�ߤ��I�6h_�k!�<p�
�XL?7�J�������u�'Y�B��WY���D�khEN�SNԶ��c>���ڹ�K`&4����a���asNn��C��k�U�[��yX��&]W��R��V޷n軡c0���u���W�0���4uMILuhŕ�>���*}j٪rM�.��(��9�[�6|�,�v7ԴQ�g��|h��b��Cd7sR=���R�yJ F/`�����WڣLp�-���f�Sr���q즤��۰ê�^?2�s��$e���Y?�<�������O�f9�N|L�"~���'$��F�����+3�����n� H�g���CU.���X�	�+B%�5V���-�@��i{�[>��qz��ٓ=}�B>�J{��1����˅������4�a���ʚ�z�m=��1�`'b��RIk˖��#��NtM��h�d`H�N��桃�C�l�4���GJjT�\�X@��Ŀ�)�ɲ�)�l}��9�#�r��w����vM���()�	n�E>��1�F��`����V��"��"�NV�����>�L=f~��ݸ�ʘ�S��2E�EL��w\C�W�<W��d�UNg��6;�LN�s0{ �I�*��{.�R��R�ɢ�N�b���O�+3��0���dGG���O5Ӽ��f/)��X���sy���S<
/�iq��kR�8���M����V���{D!��Y8Lt&;�v;�I;�/�oح3<�/z.��<�!�Y���J[�Ň�{Wͨב����>��݅9��RS��Dv��W���vL�Ԗ�d�6��U����ra�zF�������:��\�򧮵}�Q�쯠p~�" �A�����c�_ �I^(M�H�vh+����V%�}�w&w��)r�������
���Q� ���@ؤ�����z�'�\s$��{�r�9mqg�D��9��Ѣ_��▜o��9��5bN���B;���֘�k��t�M�x{��\Yr4=i��졚��040�QMĂ�jbj �ےH�\�ߏ*ƽ]��a������/���e��?uv��� R��@�[��o��wM�`k��q�~?X]0�[nu��A8Ϋ�#9W`��3��G�)-�a!D��o��~���ƾ1g�QK1�g��P>3��ϚP����!��� Lb��B?֜�J�U� G�j�\:ی����N>N#�� �Z9נ�53�jR��A��c�ͨ/����m��V0�����*����*qO�>�7��\����!b�(UT=Λ�!L��\���	B$ڔ4W��#��$���F]��R�>�4�5��3c'۹���XuRa������]��(j����g�P�j��PR�i�h#�3�N�k��~��8m��j�4�oC��?g�S2٣�Q�c�b%��ŝ����$0 �g�!���aϛ�`�s~�`@&-n��6*#\�^x;v*���j��u����<U�����ePS�k�8�RH!	��1/�r��'Ը��r�5��ҽ�T��?�f}Ԕ[����K��?���v��&�g��{2_�8|�k�Iy���~za$����ot;�PX�=0���_�7�����D#%�.��Δ��0� X�t�u�89��Нs�y�J�Hծ���!�|+�NV[��1�r���R��4��� �~��'8��+1`u�b������S���=�PC���=��ߜ�`��7��PXf�G�E}�l(.���	Xߘ�f��]�$�lVsS�$1��0�5���c�~9�@鄈N��׌�W-����������a��y�������P�$����tb���]��	"حS%���Eun�
�mC��z��e��^��v���'���V��c)�5�эUU���Rz}�2�䏔s0�h��5Yf����%S���?[�C���=�oIe�-o{��I�\��k�ʫ�A�aZJ ,�6��ڢW�R˲�5�.�v��!~��
J ��i�~�È�,��w�*N�I25u�(K䰑�i-���I���x8N��U�A���,{0Z?Q��b^�1QLiw�L��eFz�Q��Q�>�-\���d����������"�{x��a$���d���'������[�v��n���"�{�]n�q����_3Km<�P����	�[�p����(�kZ����iG���Ԯ��� ĬӃ�y�t�����[x�O �K=e��Pz��1�ϊv�F�5#�Թ�\���w&�1��Ĝn�zK�5�g�v�|{���:pW;��-ӈ<���Ѽ�̓��5��(幊(>��!�W���+C�����-ȣ�Xp��,LK%fI�
{�0�Bn2&�7����pS�U5�Y�}�r���B�.k!C�~�������d�Ym0�X�@��Ȯ=�UВ�N�*8	��I#� Og!�X+�£�8*�[G`�1��2��!&��y�_���h���"\=��7�5>�}GBt�R��g�'S�[
r�;dh21`���wu�֙��G
#��䚅��SL�YKT�>��h�p��S���GE�0GR[�	^����q�( ���ᡣ#FRQf��˯�8%UJ���a�>&�ά����]�B���O��@�{�p��-yo�+�p�M��ٛz���ў�wP$e�℞���y�=%ȽQC��q�fKf8��{C*~JM�#k�$;lǧk<�D��B/��Ħ�Ee �Y]Z4bv��s`r�)-�ޟb�@�'E����	�@�`9�5�����
�j7� �;xs���9=|��1��$
R��X��$��b�CER@�Y��
��Av��*k�2E�2��Cj�Q6y�:��Ö���l��+1JG&�j�H���D�%�ǝ����?���r�%H���3�5Z}��k�g��)y�oK�}#��i����I��y��+��4׃�{���:��nk�Ɠ���$ �>���}؟����r0��K+�^_A���4.�~�������R* ֩�v����^B2����g��' ��{�b�o��������^!��e��0�B�q������KjRJ��.;`�(�2���bb��:hJxr�X���D't�����,�_4��@�U����b�"ױPN�VT'�X"�Q$��k��0�`��,
���j�S`o*��8V����$'1'�����	���k��h?!~/3w!�C�����=5@�0٨�?~#�n�lH�= ����#��e��h,.�ZVv<���liss�F],��Yn�[��4����i}C1�f܂���,~܂k�)?��S��T��p���Z^+?g�V�o| Nl��U�6�����u|$b�ѫ��y��K��FT��Ǚ��>�������}6���1$�Yd41hƲ4V6h ��Z{�b�˙�߷��+Ҥ�_i;F��&m~b��N�5����a����ޓ@����Ӥ��K�EꗕY�Ƞfߋ�6﵈��~�n�F�y�6V~���$��Hw�	�mz�4������5���J�?y��p����^Q��X����8G���q0+��2�|�G�(���d��"h]N8�B��q�9�R�6C�.�{�ˎ�PB�Ec~?���ܒx��)�%�1�O�>�U>#	n\�E��}���Fr��)Q��ͅp%)�	���>�����	YP�z�;��+CC�&��Y����2ӟ�U��0e���u����8nJ6p>�'�!jM�@�w�_���V5�5���ßY���Z��/�g.��T$��'5���h
��y�lC���k�P�;�� ꭰ��B��ݐ��-�J�Wa�Ck������G��e�^m�]��������#L����k!#�Hu~xs�^���,�*��$����Z�!�	���
>���!�7xz�e���H<���A����g!���^��Y�]\�l���K���j�)>�I�ET��k�>����;�x��?˒<<I������T>D7FaS�Í�o��=�)q�{0D�vH;���J�X�V���Y�K�x�>y0�.W]��� G��4-��-Qdx��>g�TSYl��+)4�٠�1Y���`����>���7��!�ﾮ�Ε5�͊��X������7h2;�� ����@gH����f�1ࢆ@�?�r����l������yE��_���ē%��h���$��b]�$��п�LxS�� .'<�۞ȉr�����W�l�����MwZ�"��*2ƛ�<#�j��]Gv��X��'�9�Vs-e��;��ܷ�o���N{mQ*4vz���,�#P�Ƭ�M�6�Ayr3�!%�%�C�|;�\���~��o͔
G�������0�����4��a�"Y �6�����(H�k�p.-����|j�J� x�	��&J�̲��	B?J�^��#WXG3�E�d9�h�[�%��#�r�������i$�*�ez>�uD4ĂR��G�� N6q
?���h=}4*!)����n�{>0�}
�V�Ds�Ҕ���<��Nr�.
C�;�
!$d�k�JO�<���C_Z��Z't(���*`�h����O�~S�v_��DBbd]���9�9�_����[�#ݫ�d�wc꾗xr�9�֗����JY��|���T�\��B�|�!܌�̮<)�k�ύ�U A���H�T��4H6�8��c�뒔J2�\~�M9-��?W۾�0�^_z7�����W��M;���ߍ=s�a�~���h�b�;e�d���΅7U_���5���)���V���c	������S"bT�^��?=�,�
��?����^d|W�G�҂��1����z��'90�nx��{�� �E�u��آ��x�;�Bx2��m�jS˄�������2��\/N�lBUNm��:�y~mBxHH+��j;�B��K J4`�gC"B��c�-��?[�:��ߐ&T�t.ĐK��zʹ{ѿ#�ܮ��;�yQ�x;����[���@ё\3���e�l{@p��I��S�rВ�:��9�7_�)�劓����QC�Y�����6�m�b���Ӌf5. �>��s��ʲ7�C�� T���梟��*p��d3ߚ&�="��iڦq������uܾe��2�Q�$����oO$�8�S��}w=�� �*�^�(�HkLȓz"F����!��_��K�4A-{gY��s�'F
Ar�@��0��l�O7Ba��/�d�nX��5�u��b�dlziZF��ᴗ����ˇ�¼��s3��D�tR��*��U��η���H+��~"�0�F˴���#w��u�T�sJ=a�԰�H��V�d���Qf8�|X*p� i�X���2�^QH��T((�����'e(������xᲥ祺+�k�[���-����oC�w�
VB���fb��Qt�36�U�,���~�<fy����/HeP��v��5b}W�H�ElQ������gIP��(
\L��������n�
�i@~��x�N),4�7擲��,�(�y�X�����9��sp�"�g5"Z8.�3f�N�4~6a�{ƉSowa�����N��h<,<a�[�:��ds�zx�}-p
�X�.��L>xS����VM�-�Ө�|y��J��E]
~*�k_67a��<�P)��`�T#o�.��/�wo�'}v-�cJu)����]H%��z�&R���!�[���C���3��7mD6��z��B�WN���5����{VǴY��Hn��߸�~0c���K��@<}�H���R�R�~��ņ�%4C�x�#`���@IX�p��'�0~^$��3�W����d$n�G�Ph�*��P��¹����lQ3/$�7�d�wI��'s�,��g6�q������rVx��J�3�W_$�cC�~����F*�
�Z�OQ��K��
��ᢪ���[X)�k�j��o%�1����LyB��B�N��x.ح���2�Qȝ"Aբ%��B�+N!�����8_Y����n|k��* 즷�o�uQTj���`��*TmS��OJYa*w]�����AKz��Ӆ�,c G,�y�h=��w �c"���޺��$G���ϐS�iLa��⓵��"2�9�S�@����~�|�GYd��^!�T�w&s�D�9����@wt�܈�F���@��;����O��B� y�eS:"�����~z�8��4U���d̕xE��c�:%�=�	�Gi���P>xJs�\�(0�O�V���gL?����z��e+�(���LUj��5�.��Md�B}�a�ot�=%;�Xƚ��^T���O�Ѥ����o����a%&R�P�`_}x�;���Cn�,�?YN�i77�&�t� ©�=4��Ç\VԼ��S�z��/�O<���B�����sgȻ�g���a,����������$MzB����"(�^Px�	�ҹ}��L�*�~&���).V��>�ݼ��B�ɽ@�$�h��:Ք9	��w�O��_��!��[9I�5a��-�j���(\�P>0)�x�����T�^����QlC�{�h��̇��.\}����q�� �y��t���ڜV5�C��o%�Y�wC*�	�Ү ���X!gOQ��hsN�=�
S[��2t��_[l:��u�{����F�}Ns�8�cæ��fz�ˑ��#���M��˽�Qo,����=�o��{5E[�m	j��pW*t�g)��+�E���)y��cJ�b,�=?K)S�Z���n�Q����Bk5��6���H:�S�� +UN�hp]O[2�^�h�eRlf��l/�����^(׮����*��sC �������BV^�����ѿ�|8��AK5̰g�tr�x�(V��a�?�)�. hbyV/쉾Ү���k��|}�Q<�%W#D��ऍ4�c�VR15���]t�_	���f�qӜ!�}X�\�6�D@D�HA�1�quU�q94Ȓ���g_���.��sq���g���ċxw�-�3��qRp�_�����AA&k��sr���ǻM/V�R�����F��gq1q(�k��6�T�=$��� y�����5��9��*J[��`
8?�%�תީZ}����R\U	�g�����0%�p���y�ڼl�d	O��sh�d��˅��$��,q��yFq�p���*\
 ����ÈG'J ��6�2�[V��ۜ��#��R���ύ�95��z����N>����ʓW.ȼq&��`�R���H"2������W,�����SVVv�&�H�@�Sb������jCd�x�8�C����܁$&���y����Y۝*�$��f��%�T��(d<I�)&�{���R�����7r��H t8'!��@'��Z�*����WLMC�"�M>C�C��6�����:|?8���K���6������D�q�ezuGU�f/�鵇�f�`���	��{���]�cY�z��-��{ s��Ʈ�х� �������|d�H�R��������M���'�{�G��#�=��U �� ['��q��^ɸ�V�������& ��kl���Ѣ��qU�A�	
�
�D���P`9�L�$\67��$���M�˨��&	H$��1���ᕜ�%}��>�{��!������`aQ���kW,V�3ⲹ����g�����ֱ��O���Qj#{졵r�wQ��VWp[6�5�����B>4O����d�A�ãթg9��h.�G�V�e�Qw���!"��mz��"�L��\q-�U��K�xU�W%�l����@s������s�cЄ(t�]�W ����?����W[���żVXxo�'��w�\�_�?�t�^A����s������yz4zA��4�m�85h*�^	9�֟�f��B��~�|�+�����ӵ ���t��4ڙ�b�.�(��F����FZ��^�.��ZR�3���)�yv������������tٛ�>�\��U]SA���Bi&s�/�(u��<bG���.�-����*���~Gx�y�oue|�j�!�=��=��9�БZB��J��g�3V��&0 �����������/!{"f��k��4�����l�TwL-c���.���="��s �fc����e�|z^�ͷD٦��[}�����CDrHW��=�#;�#1���R.S��)!oQI�̔��'z���W��Y�[�6���?k��&H��u4� _�G��V:z]�}��tV�G	�z��`6�A~|n'�Ouz�;7���U�F�����l���#~�Xvb
���&��H.������-����zQ*EBC����/[� ��"L'�ޠ�y]�{���:��sg����	'h�u�DM���`N�f�N緌�U%�[��M��7�ris����T(kh����w�[���t�Cd�붘#[9bf�s�F�Is�:1v���ÇRk(P.b��?<S�p�k~�B}�FjD���n���,�+Y��-���#��gy;E�S��`}��Pd�û�S��\Y�&m%֬���	�/z�:�fR�]�Rg�b�4R����-��{��$�^TӿfU�w�R�1;��x&s&A�q�X�C�A����;���B3m�#�d{���d~F�ʐkQ��op���.*jξ��J����Nv���y�f�N����"�.�˭>�pI%��!�ua�J׉Q�,i�UA����t�.�����%��U4PM���i�P?/bXq����HI jݎ�����䠬C;���f*e����	C�S��,���g�*����5T�����`��LU)���K��tO�Phf�����RZLh��23�3�t�4N:����:�(E�Jr5���m0g�FS������+�\������rl9n<�n�\��( ��,d�����k�장�u�i8T�����쭔�� K��AI�t�z�zx%�%z %S�27�/���k�ʊ��XgP�N�y��Z]�R@A�WZ�3�?�/�m����d�]z�� ���\0n�Y��Fo1t\D;e,��%�q���h�	UO�Ȥ�Gr�'���aǾx��ʟ������gctϪ1q��f����"��B�X����
�����Br�^��)6��C��a$\U&��O���yBz���_�0���L��Z?��	Z�(�*����Cw��*p�8��%�f�,��L,jq�`
����g���<�(��U�����GfT(&A OR �D#x��%61d��8dʀ�?m�*�R�-�ӝgzu��'z-���V�/���tY�T��F:���gtP�U�XAd2�,��%psRQ ��'}fO�Z q�K��"��Y�ݳ�
�g;"���Y�}Gָ�'I t��է���+�N����1de>�d�Z��nf����d�[B�������5#U����j�WO��B��>�[}HXY�U�[qf��`R�zsj#l�Vc�s$B�;�aHֽ�����ơ�b%bHؖ�<�^V�7��@�F�5i��2w��/�D"�٣�;�򨃵ZI�������E ��kG�c5�gՎ�q�����(Иq��L�0�&z��f
�	Wp?�SJI�:����I���OOr0}tV�	����}Z�k������[AI����V#���P�7�8�_F��d���`u6M:�I��-$��Gp~��fL{NH�=��L4����Q6Kx2���G�g�Ճii�.�F�S]�!7���Z��I��W�y0�M�Z+ۛ�K�
��h�[�s]����"�K�c�k�7�`6i48ڵ�z���&q�o�9�u0�Ƕ�U�W.�4@յ�6\O,BR�(�e��·h�i�g)�����b����0P������x�DA���7z��B�=�1�$�:�M̧F���ã��A�iI�Y�ҿ�hh�v�F�#��Z�2�}�z���Aݒ� :��fM<Jjۧ�`�ǅ�H}��s�xڦ�4H}���(ܰ�A
�;����oJ���Z��!슮qە_w��X?���ڄ� ��ʠH����c�C��,�]$��1��<#�l�����:�ٚ�3b�xؐS��"�X���Tq�a���7ӿ5G�L �G��V��`��E�l�i�T��H*��$`�sG��Ř���\����� R±�(ț��|q��j-�D�ƍz5t�ט7�H0$�Wy~���G5��7�q����<g0��7����~�N�Gd��
�Y���j] P/�36m�e�dW�cۘ�W���b6�5�_芒y�r	���GBq�r�6J`W��bks�a+!�Xl^f�5 �6e� �aI�s�Nr(�g�3!�`���4(�Y�#���剺�k�Z5�g�w�"�k���b1'[���T��]�3q����:2Q�PM����c�.o�|k;��Di���$�(�c�I�;�����]�h���E�g8�N[�*�Ɔj�^�l��ȳ�<���JT8����'44E�P��\��4+Y�IJ�DM 9gz�W9�<G(f�5��N1{���/��Ћ�.VUH�:�Aېq�e��!��~�n�:RZl��v�}��]\	�k+5\��9Q�k�����Y�nk&$�Ś���Օ�ו.��������k5/�u
%����t�$�$��͇6cI6��1b7�f}t�~.���m�Z��I���3�Xc�����E����4�.��dzV�=hu��ž4�刼k��>�fH̳kq���9)eIq���O�>Z\�5J�7%"֝�m�J�ƒ,�m��"�]͎J� ��~l�P�<,�U���b0�o4(9׷�o}�Ôr�.�¥��M��]׽b�S���S�F�����Qi��_�U�������c#+n��c]Q�)KZ͞i��AD|b���la���c�+r�_���Ѻh�d�$�d#�o֦Q�׫��p	P���?�L���`�]����;l=!j(�Q���^��-B����J�.b�uH
m���5%������-��Zb4�?�*��ա|��|0j�F�4$J�[L�Q�v!|���ʓ�<M���?&a4��I��Y���e8��2����5����~��"���~:]T�Ζ��3*�:r笎H����ƍ�|�d�~���E��}�?\��o˦����������Qdg��lrE�O^�H��o�<8���r�x/.�>�0,���3���-�]�$ޫ��H� ���"ž+.��"(G���}�a���qԼ��Mv=g��3������y��% �	]���gj��xA�T�$�:L�]�L'���i:ێ����h�Π�S|�%xɒ_;s���rٜ'������k�y]d��`�+��ɝ�E����i�2�w(��U�E��������'@7<9Y)��O�n�AAu ������DP8���ӊ=@n'�|�,DKV�%�~�(�8�]��W5���;�a���4��O/� ;��n���$:1~�x�<��s@H���GnD�l�P���!�K5�I�533}h�,4D��f�N��� ��1SNMd��Ck?�W$t]oL3�圤��n͝�B�����D����r!�M��)�0-.:@v\�kV/�l�k�ׄy���8�+\��+(Ȍ.������_�rz۴i��I�Ӥ�� '��?R��)n���Tr�I����ęE�L�֯9�q���sA�T�3uV�!�"J�!d�� �׭~����������B�^��휄Y
� ���O��N�מ� ��N��Zȧ�� ����Ļ��;5���m-���[� ,Z>eݜ������?�^���%�`ʌ�fܐ���-O�v���3���~�;��]�l}�!:Oy��q4�c��=���e̛>U1�a���K�U�*�| ���g:f6Ƥ�q퓩�H�'ڄ־s�[aʝP�(���%He�C��B|���iEWӟ'JT���n�!I����q�X�US���6����)B��Ƥ���	��2������_�S-(DJSZ��"iu���������)d�d����|E@��VIk�����J���E~�l�������	��\y��%�~I��!����k��yΟ����㜭&DY�:��8��{��w�^6��d����F�l'�#���i��`��7�#�@��6�E��'��o�'�o&��N�E[���e��*#�[Q�	��|nƾ"�ʈ,A�0�����|�[����8�#b@�^0��N�'c!��)$��D����LQz-#�ظ��1�oPŘ00�c��t�$r*�Ž9���W9ۄ%��ٜ�7�w��1w�-�#��^Ѝ���;�kg��� �=��"l�v�m�rހ�B�!*��1k�y�G7�+[��6�w��+R�m5����Q�T��D�/?���ǋPld�m!|c�i��K���'GkfkaZ������l[UD:}s��I�zV�L����:fܛ5x�ug�M�;��Iƺ=��#���0n�����[,��t!��LTA5hW1����.��x�U��xޗ�>��4���7u�W]W*�M�V�R���]����zEc��'��j�$5��TX�5��'h���tj`�PVA �m�)t���r�r���
��'T ��#s��X��� iO�͠혊h�U㸤����c��s��.F_�Mrf�_���^��wkP�+���o��C�R+Y���0�r�v5p6���s=��������[�z�"2�%��A��s�qN��*��М\���*�.'��>��n���Ua�%2����Yb:6��ck�����e�)В�=Bu|�����k�?�E�]*	>٢�9���\$ZU]�> 5�!�|�z�#CP�5���Z����>��M���ך(�Nɭ��V##�O������@�P~�X߿�����<�cO"�,�V����¡�i�X<YQG(Ǒ�<k���l snX�Al��u^��T&(�J^e���Ec��k4�/Z��n��,<#������0�����A<ƞ-�2�zD3���*D2�)Py��k-�{vK��6NHk���W��'˰��]�F.��M��4��Ŕ�x@g�)����t��t�;S*��2;��N�x'�����h~�th�b���-Hy�aJ����<?vM��:�B\ˎJ���t�1
{e3����䥆��d���Bg���T��)y�E�dp��@5o�!��r��L�[
�ˀ���+su��9TtIUD��w�R�q9�A�����g�^{mq���ֳC����=�>�]и*�M��6��r�<���H��p��pP\#S�f��Y�Ү%B��FY�Q�q�$�J�p\ɼɴxK�o	�WM�M$�ꉖh�2&�G|����+ s� �8�ۧF�\�������e�U������3'�H_zԸՆ�Of�G�mw�qDxY��,�y������"."�Gͫ�w�������h�M��q\�$m�s��7D|�I�v��p�'%�����l��HlL�𤒪�E���A���&Zp�⦅C/��b.GD0N�:z2��@bh�Y!Υ� �d3K�!�����䛠�Ko�$QћM`_��u��=[6�I�\ズSw~��8���-���F<u�<����x�޺ـ! '���]��̂�DJʌn���n3<0�L(.��B�O6���� EDǤ�����+��+���x.�|Gh�� 9���'���ؒh�P�B#�����	����5w��]!��$O󞫉a�l��r�����f�1svEo����8�^��Z:���ܬq���S�LH��CF�9�`�R�a�Ȱz?�\?F̍b���fTA�=��)f�o���G �����˄� !�*�7�%� S��Gk��� k}lh��#A��W��*��;�
������95SNv	��R�lΫ �d�I���L8o���Z�4s�M�����MR�v�)�3H�����H�q�i�=!=֡�x�g)�e d����I��������P^(��B���+���-��\N�zqJ;a��t�$ް�l��s����hr$�O��tD'Z�U�����ɐ꽉m0G�155�ⶍ$�J8�:f��l}*�o?y�,�A��X�X��'lJ��H y�=�R5K0屻�+��)Zfl֔S<�ߐ)�Bh���S_4�&z\�}n��yY��3�(�}z7�l�J��X�g0�]�:� L�y��4i&��.���tw$�eR�&��(x/(�6��Q�hF�]Gi(��K�\��P��&�5��ݨ������y.0Y	��e�)��&�|�^�Y!��ֹ9� ��ZN����9��/]^X�R������*k���p����Aߚ잍J�ZH�)H��M�NU�U�m���ܭB�y�Ҫq2y��@��3}��~@GeS��$�ɰ��8�*�"����ӮW#�p�����f��%W������3$�5lL��.�vJ��7��Mߣ=�5�A���Z�0�8|�YK��5;���+�����[Q�R�L�Ѷ�����,�mZ�Dr�FB����R��-Ƚb/J2ƥlۼa�L�ܹ�PmD{K?d���DL�-�5�kH � >�9���K6>�D�a&�K*J��~���es&�/K��X��^Y<�s�N%���+��w�0�7;���v9��̹N�A�?F����������qU�p{�V��N��� AʈK��Uw�ؙ��y��Q�=q�,0�vو�I�4Gl�wq�9��6��/���K���K�y�C�գ��/��a�]�^�.�ٹt:U�J̇�&Vl�}8�{R�e'��y�of�Xt�Y3�z��zqs|9�|�p��� �ܯِs���9'@��2��_f�?��}�Ɵ�� o�.�y��>�,y�����?�N��K���F��6�3Y�dh9t'��uX�;�a�N*>�P|i6�@d�R�$Q�8�!��NT:+U^�yƄ,���R�`x;�����1��k�����;����z�	� zn��"���>�c��a�7���?�v�`��ڻċ�d���K~tSI&lك���#�Z�Hj'^��A0Ҙ8gh������cЂ����rX�ȃ�彰:�-p+W,���� �eЌ�f����f|��"\E�8��B������xY;�YR.L���!�e�M<ޚ)ͭ��pn�T�I\C�5n���:��E	oMSrp*ڵ+�*����ԓ�����)�0��/��"i3y��7��1��b���2�ryC�@4�=v�Z<��:�j��aQh���"��
��9&��W�;����S0�ܫE��,�8It�-L�O������(��E�չ�7C�h�TkN�רYȤ��h�wW��(oOŴ
~WZ̙X�ԕ��_��U>#����}㸓$_��d녺[RU ��m����M���N�u�l]�b���`zJ�M=��1�����-�Di45��0�� S�8s�}�2�5CW�;���p�Q'ʼ� ˢ$����B��ݚ�J���uc�k���|y>�4�/�4,���=�>�= ��g��b�ܝ��
��r\;�RC��*�0�7��b.�د��rVq�_�VlU&�N�n�Μ29�_�����|9�*��W4��W��JيY��5�-�=�j[!E�0��c��L�U_|OIB�a���4$�hC��&@i�e��I����9�g� x k�n�'Vs�ky�M���+ɬ�ґ&8Fs���,��#%���DH��޴��v�1����:�n�?����7L�p��_�7A�Oޑ�Q� P���y($�-!V��r�a�[�P�ؾV�'���#q�Sڻ��-�ۀ�����B�s��)�(z����,��9t	���9h��q�6_���-� sX��l����ұ �u^Da�r+���ct��o�>�0��PL�w���ׂ���D�3>�A	o��6�`�I��z��	N�3ر�n���36­Bhu:�a�ȁ+B��0ԩ7�8��\��`g�O=�mpӴ���D��r�N�p��A)<9-��|{N��[Gp�V��2�B�"jFS�p�� C��&��ŇAS��2�:���E�*6�	�Pş�����N_z�� �A�p�ȑ��~p;a��]� ���A��g�-"l�v��1�2���1^ˡ�Jy���`
����2{�X�
B��!9�YR�`�����|�<���!���1�k�9ɘ�Sp�	�ʼ;�UY�]��	J�������5�����2i�y'�RKm�:��#�t��ٖ|�>�q��o�Ͱ���������.�B!&O��jQT1T�7���JD�D���}g��|f����9�{���}�����w�ܧ���Y��K''���`�MWTAE�L9laۋ�(�Xw�<8r��N�Z5�X\e��dg�����;��)���u
K)R4�7uT�$�چT��$�F�,#Vl�>���Z8��H�跎ܖ-.��c�i�o,���K�#?��?꒢|hP�3x���T��U�S�-�Ȳ��B:��[����¨�l���&����.?~����f�a�1]xKY/�� �T|�����Ky�'>&������:���Z��M�`�+4\��ޢ�*�4S�Ȥ<�Xckd����I�@̥��L�ф���<�z�4-��kB�hs�2=���;�		�x�� 	�{݌@���:;��>�++��\D��5j�#�S�Me/v��}����t�������Д���$-�����}�hkRW�5x=Fj9�Ұ_���l>�^���u�R����m� /�h�cgZqy
��o�����ƶ?,e(]���>4䨌���q+*�)�9���{�<���U�,�H�g���p�-W�ͣ��q)y���l���P� �	P6(���zd�Cۭdw��<y��&9*�~��_��s�)q�5�Gx`(puV��'XPI��(�����#��f��K�$~z�i���.�� M�n$��4`�ζ�˨J�۟퀆������"��b0���1�:7:��KÂh�b�3ϣ4d��ځч/��������ɀs!�OP�8���?����K�(� @5#K4ȎN�,��4av�!��(��&,i�S�n�e�W�f��U�m�F#��[)!&�Ƥ��[�1^eL���Z6h��dSj[㼾�u=�yVD���et?����$�.�Du�k�f�%1:�hB�W�麮��-�EWcf�����u����kT����L��o/>���h�C��S���1���p�j�+9���/0�|	���B�n�1W���r	|ƒ�X�(���Ҙ����|��\�eu���T��Z�6-�j�L����ă�p�P$yD����6�������c��K�D� ���7L�)J�)�"_I\ѭ�����̠���Xs��d�"*����=L�ژ�il���@j��*�O6�T쳪����ՙD��8ᘄ�?�F=��)�*a>s�3!v���͓�-���4B�,[����E�`(����Q]�cG�qM#+�������g7$���[n�H�X �v��� /�o�i��!���Oa����u�������2���<�� �+z�F�\/Ы܄rN�Zf�q�hPh`�����RA�
�J����n�ޤg�.f޼�Byל�^r�W<�.z�S<�)��ROA��Yt,;�L�Y�4��<r���P�TA9nHĵ_Z��m�q�|��Oz7J�1��!�����?*\� �.1���N"8�a���;��W�����}<qq 8��9ux�U���pB΍�Ɯ�Z]��i�;�ї`	�k���g|�Q
[��+��{�P4ݷ�4 +�m=^��2:��>�o/t���ڣ�Чe��BdDt�q����
+1mlR��m8�e�[���R����dS(7��D�)fX�o��7��4��j���s-��[�\�i��J�����I��m�۶��D�Ή�����fc���Y�����i�tV�
��ki%C�sC��'��,۽��
��u�e�F�7)k����-���9B.B��XI��H~�ě�����mi<~,�_� ��
���C�ㄐ����D{8a���R[�7�D1�eA����)� �
Br\'ȿ�"�Y�|rs�"/p�2
P+�SR0�Jyp6q���.��f�B��Ê���GW����p����e9������ y��R
5��ww�ˆ,�A=��{4�N�����}������t5�����7��:�ަ�W)�	� J$}�/���{/�y�l|/��	[ʅJE��a���f��ΖI�>3�	nr�"9�v�W�y�g]��Į�'a.Ts^'��9��bU���EU��Ji�?���T�J��>G�N� �fpݼ_/O�j�SSxx�+i��o�\�G�l�gݯfЙ��J��Z|�E�^���H�]��7�
�6�����>�r��c վED �S�D�/�N����J���إTB�/�g�����ה�Zթ�H�����=_��,� �t��O���o?8���;.g�����}GmJh�ʦv�@	�r�g((=ە&&��:��>_/��
�62P�I�g?�c�@� ��t�	�-�-8��p��Ӣb�߶[�^��}2Ft���\�)��"���>n?�ԓ�b���[�`0C(����_�%T[���"�ހ,�[٠��:hg���E��q��2�1 z��A�oTu���J���Ph��t�D�>`Z�a�`�y�\��O҅I ��.�2��v��/�R��y��J���h����蝉8� æn�9���ݺ�p��%��02`x���"&0J��!�4-$��Օ��e���R���b'��nf;��'��8s-��l�Zū�z� ڬ\k���%��̸�^r����W;'�%��0����=/�d���6�+�I��q:��$>�zx���ʘl4Jtݧ�]��u�|�#ŏ2�]m���t5�@!$�@	I�#P�Y�����)1�&�;�H:.����?W �m��apt���x�,��Bjy����c>29��ǘb(a{�U/�g�1�'�þEt���^j SL(a�ϳ��:O������_���i,��h�T��#�]����5}jl�d�g{� k�E�h�� �w����P�S�e��ALs�9�v�snj�N�#a�&��\H��p_��,@�N�<��J�ˬ���rK�z�QA2,�eTh03�M�RȂj<��:&4�9~�/���<��d�'��7#n������ɹ4{���F�W��ϝ�ǃ�%��&��s7����7�J���db��}��*Y�J��6��ϩT�+�[�>��w��"ҍ[��
8`�pa�Ϯ�SB��� L�����9ԄL[׼�1#��X��^����y�2էp��&�j�o9 ����UpE�y��ٗ����įMհZ�k��¼9i�(�V��
M��%!�f_l�e9�O0l�ٛ��V�A���ŕ����U�fk��yh�_�lE3�$@��W�� 4R�)�a�/y�����.-R�]3�̰�y�T���>q���?+O���)�w�22m\�b'zZw@�a�+	��i��_��-�"�s4V�Ak$�fO��rj����e�S�SX��=:�/�9��ᜁrW��v^#}�[nzr/ֲ����O�ķ8❬].@���;Y���a}�\_���M�Ap9gG��I�:$zθ;��r���q;��爟�����<�tܜo����T�V�H�ƍ{��
$y�����>&7K��K?B:*H���5w��!{��_���Y�(@ó�rp��|^Lwx�bU�H��:�Qi^���Gl�ُ�dc��V���tx[��Ы�^�?0���׎tIJz�G~��xjd��G�h�������%�Z'`F�2o���*����k �b|��#轭���D+�%,�i,�b$�؀ �����N3�dʹ��}΄Fh�4��RE�G���s��b��������3y��Mb]Cm�+TL���'H������;!��ke(��巾�ȵ�m}�;�#;X|���&T��/_s޶�����?=�k��r�1�0�v�Dm���(���$��
=�K�MF�x����O	Lۍ���h��?.E(L� tU"�F��	��j^x
�I��)P�1��q:WF����mu���{~�$�ӂ>w�^�5�Z�W���C�C�i:9Au���!Өo��8�Fg���f8�Й�:����Q�u[��_ЮLU����w�ɿܜ�{|�V`�%����*n�${t��V�n���Y�t���O�Y[�1$�����'�|:��Lj��$��>x�V��w)	rJ�J�$GIP����M��p��a�3k��bSL��6u�!$�"o�AB�4�ȝ! �P���CH�\�.�h:����v���.Gvl�E�,��)�o|��}\�D��	zz��6U�kS����'�5Q�'0�����YhqP:��� $�-w��R��c�("<�ذ������$�X[�&W����
�<��:!0�����-cV>�f���s�ʭ�4+�K���>���{�~&gi:�s�#����C�J�ȵs��]f[����Z溇����;�Nl>��X�#J��v�� �5i)�$��Q�5�Wz^x����t3r���T����3�ԝ�1��
���k�wA�!���6��y�Ak�`�p?����{0�R8O~}$Ty{�KQ���'���ܗ[sp�g��	A!�
�!�˫=�U=�{�E�,l�j���Ke���"z����Wğ��F�P�g�d?�$��:@muU�+_r��Ǆ�q������V� ��}v�G;[�KM��;ɐ��#��� V��U׆(#�e!�H����h�<�c�o�E�5Ay�ј�:��+<�`��[=35�c��c `��(��H�~���񫌣{
�{�����ʡ������aS��j��IV�v�l �LNj�$�o�����~�g;,��D�]ۯ���菱
��ٔE#�E��m/B�*��>�g��?�/�l�>gO�g= ��+�@��<�v�V�D0�px�=/������m��*[�2��w6(��d�.:˶FBdY���]r�n+�h��qh	��o<r�{p��9S���u@��������:Vb_Kūr�z?Sřf*��AL3��ʌ�>�_{��ۉG���5@��fn�b����t�[X����vl]���ufuGe�� 9Tl��M�E��p4r�8��K���0k���o��Jb��4�|`������P�O� ϨM�/V ��b5�����iP��8�=4e����)B�Th�30�Q�;��6������$-?��8�\�joٱ�D�j�X�ۻ��Й�A��T����������"GN�*a�CLj�W�� y��)��#&���Mt˃��	kJ���%����k��ʉU�þM��t���X&�0�p�*���Ҳ;`e�C�DF�����;�'f?J�>���ƒ�#�w�ƾ7M�s�B1Q)�)>���v�D%^��x7�Q�+�U���ڡ�j�msvh8]�wv�2C�-� ��؁�/�6����K2f�0�2�	����q3�[����\���P���@9X%2�Wr_�<[>�?^�{=0D�y��R�̉�bg���a�4y����Ws�e�L�2�N�-�oD�Y������cHd1�E���&���X��o�ྨd�&OlŻ����HK��|��\-W2��N�N2�7�)�9��v6^-ݹ!X7ʃ�\�I���o���K$��,EQ��g�t%٪�d�ߨ=q-^�a���U�����}I^��>��:I�'ˎJd��[��r��IY�%m������������P����6�߳ ����x���¢�����|>L��� ���W�cŵ�C�HF~q��%'���9�\�%�C�t��xM#ʌA�J�9|r�a���ݫ�v��W&`���(�\�����D��k��+��b�����q�Y���"��ry����p�;�V�.t�-
��B^8������c��6�k3�0�]�\�uPt/h��{#[w����C�5�W�x������C!N�r0=��jL�4�����X��M��1}���}u(-�A�,��-�{;s{!Z��B5�qL_/ S??�:|�a���K씹���#�z�|�kQ�sy��u8^ �N�u{� g,m'2����~�I.)��
�J<�վ�R�HǓ���D�p�
�Y���,E�P�P����h�U�CF(�nⁿ�|��Hp��u^�6���%��+����X�Nk��5��@�&���4�5ܪ���2'��,�%'�2e4�� 6!���[�V�]
�/�Z��Qv|yI����T㏀csy!q��]�֥w�4�LnO�!^���me)�����D��o���`h;:�ĩJ&���1`=�D2�oNz3�ހ�+`G]�{υ�q���,� �MR���2A�g�E�������D�immo�{�L,S��OT"�v�!ҭ��NOz�įV3��Ц`+s�we$�p�^����F�C[h�
�^[劘p�㵬�ӷ�,>P�e�SaM��lp���2w)��m�R�n�0���9p�9�a�9a����4�%���(��e�T�{���6�|tcSc�a\w|��G��49��p������<隢撘$a��t�+WN���L�� ���λX0�	�o�^oK�S �Wu}�f�HV^�նKtUI,�X�a�����[� !�Ɗ����8OFDYIy���`R�GF���8���rU�}~W�b
ԶF�.+���%�
�9�u?�0~j�����M�o���HP�M�TQ@%��h���8�'�B�Y �J��T���0Wj]�'J�Q��_��S>���N�l�ѦTvc���v��\LuVd�@��<|Oe���@���S�Svd�+���1�Ԭ�ޫ���{�1/B턜�y�S��b��!uR�4��Z0����EӒ�:��~j�N�88�/�D2�K೛��{�Q�WQ��}C�s�?�=a9�xnH�#��j�;ɇH^J�p6o7.s_	Ô+�*C��p3d�Kt�(&�Qɑ���W!��;��T ��.��u��pW(�ny'ee.��a�^�N��k�l�L��(%�pG���9;�)��z���U-���W�o�T5��GK%��P2�iZ����%Վ���o��q�D�S�-�O�s'%�3�r���ژh��t�vD{zU|�q�����g	��wG+`�1��)�`���!�Y�bp�+����ͤf)O���>ƁtUZ-����p��&V�/��2˝��m	�<��ON�H`�����T���[���w0i�3�K��ߩ{�!��|�B��B=\��%=a�4����	f5�1	"pՓ0TY	��C�j�9B*wv��8z=��؜�q���^�|i��&j��=`<�0�Ե�^~<
�]m��~�8�]������r����Y�"kw0��oi��	ҹ�Q
7����C:.����/�v��q�+u����v�D�9���ᓘ�m��ך%�EQ{�S*�2��Lx/��D���D���wx���s8!v��r�.���4_e��@V��U�
e��5J(�����^����mv����=js>�4������S�+Ĥx$:�˪�@�}lq��ћsP�ݏ+�e�X�e�ʡ��^�a$@��>X�`�Q/��\�E�C�K��b�������ȫ�e�c�)t�!�AoS(�P�k��� �4��Te{���{��F8w�k��B�Nr�j����/��}� f�y�v���!@L�gc��_	��2��d��%�cG�?#�w]�h#m	ŊN]{��()��!��Ml|+5l2���"v��c@���<4SY���H=.�K#����F�OO^��ư
�{�4K�Nʾ%\�Ɯ�ޡ�l���f�8U��}���y�����Φ*�}5Ǯ�E�rt��Ɗ��{�f��9'�"�{�F�wھ����>�W���& �l ��Iu���FnGM�aTN�h�WX�
|K_t0dԦ ��O���X��x��m��}���!�tɓ��;�p�i1�Pł�k=WK��3�F��^�r�펄tH�M@�!i��m�t#�g�u=�x��Gw'a��@SM�>�.�k�>��Sa�P���u#�s�c�tޥ�P�j������g	���f�!N�q��[�'�b��h�m��T�SW�R��W	�W�� ¦�ymT�����2[�%W�lk{v�j������|�=�8�"`�n�t��Q)����UOT��	�ٹ񎕄.#RK�i��
���]�a���W�85�ꦿ1�/�p��<��W�w�`�M�FIV�_jTSS��b�#_�b���g�7~Bkhz�L�h#wEKC9�����U�Sz�Y(��l B�و��"��QҮ4�����+��K���8�EU{q����C�X�C3�t�����OE1��v�hL=�ٸB�^D������I�Il�0�� �k�٤2���M��9tۧKD\ַ1t����!�VŶ�m95p�6 &e��NcA�.W�)�/��Qw_@i���\Өvl������:w JW{��ٌŷU8*5�V��(p�`�Ǜ�[	��Y������Р��MCq�Y��!��Z��4�����T#O�k�I\��IX��~��
�q�П��h_����9h~|�%�儝�$P�ɨP�^��l�;���F��b+T�bR��@��a6��əB#�8�H�E3��Lԫ،�O�ウ�ɹ�f�
��擐�e�fφp��K��JA@��vj1��'(-JN3��D�_Ix�2�ď��%�!L��VWEp�p���iS���լ��(�&��U�^"� �"�lv�~�FT����n|fP�xn nT'P_P���
j��Gf��I@_P,�Ws��|�����v�s_��9��O��*����:8����#��[�}{�3�	���MZi|���X�7�0{t��a����v�5Ѭ���`�om߹+	���>[Z��Ȑ�(u��$A���_�jZ�����;�@9/����ŇH�?�.F!�������Bӗ� �֧{�i{t��g�F���2���$�rW�Rjx}��c�˓���Y���T���OUO#?�a81s p|c��V`��p[�G��O
�`n5
;�,��:�_��o�Y��܁�7*~��Q�W!U,e�
:���b��[5�Ha���dy��	g�e�1u�M��l�<rz��q.q0ut��"tbd�J9�VL���5:�Ҭ�������b���]А�f�Gsv,Ñ�!Q�z	��̴QuGg�?�}E�H�F�E�6�h}E'ϖG��Id#�Y���M�Nvȶy�ñY��
��G.e6�7��W�iG�"���vE�gmJvD��.8��5K���R��|s�r?JF�+����$A�����������\���ފ�(���A;��L�i �i�̫��ay���7��lK��ξ��q)ڭ�*�/ɖ��mF�#��ً�}�����?WE�'���*sV���+���O�
>�����~�1U@��ﵐ.ă�d ��I�g`�q�b���|��%A#0�&���n�i<�>Z�,[�6���I��WC���
�(��Ӄ�<߄��J�$���o��"q(�����^��3\�[�_e�����M*9r��S/�y[z��К/<w Ii��
��D֫4������_�B���Y�@�e�ubD����F����J���)�|������M*OPk�V�L����"���h�(��tg�M������ ��=���h�E+�11�i\�e��a$�}	��v(Z�2][z�q�]�i�����+'\�Z�F<d9��*�ʈ�P�O��|MѼ�o��P=�����(�w-|�-�h��M���M�|��!�x�v�A��wS��>�:���6{�D|�s���8;l��#��/Y(����'�-. Ϩ=9�-��'��8H|���x�p�y�H��cj��h#�t��cd��Q��z!O7�Y��H'IBF��6��� B�	�=����k�8�����4�6���^�(db��2lm��k��&�ڲW���#;ؑ V��G�����پ���k�����P��{�����A��������od�\2�c��������Oc��B��P&")�k@��W0�F���y�N$5��]��"{@�	7Q����>?7u�g����%��+�D�P���q~v��L�juy��|�\#���x�ߚp����
kw��hV��9`�3�"�JFx�zy�1Z��(���W���d��X�srX/X�^U����=Fl��a�s]z��a�3>�F¹Rh���Y�3)[\���Z?a�;v ���新ʙ�MR�|e��%�������F2ix�jÿ��T׉��v��������k*8|O3J�p����L%�f�Le�N���ǫ~N�bv����\N��M��١�����$�|�'$-��5Rn�Ij����c�N�;{�p�ŧ�4>D|��.cAb�l �ѽ��P��)�����٦r`Ф�)��[��������S��_��i�,	��(���8�;��J aC&����+�H4B�K��D�Ł�J�%;�}ɕp0)��6�s��D0X:Ga���H�m��/� $z��RYN����Smڷ3���m� ����ʑ��7��2i+]*���3�{;a\����|�컬�*�$�|��srGje4��
���_�pO���o<��SX���Ա=�
�WS�2l\�.,�ҳo2*�w_�䒕����kK����5�n	�v�x?;�,oyD��+��ҏcc��1��}6�{AJ?��4s��E��t��O��p�Ⱥ���|�'����7����.��h�&�Qp�C��r�h�>��l0^�����]�w�6�K�2������.!&��㊻C�s�����sDZ����4"�s���ɑ��i��w�|�\����@|��I��RꮝG����3��)�;Ch9���it���I@(��4�4	��7}�Q���<�;�����7���$�!�vN�c�����t1	�����������\�F��Ӕ/�E�Q'����\��J:sVB�͞a|�!�i~͏���*
��8��%EdZԡ�u+kT���~�p[�
��>�T��t���x����ϔ�V*�X�[Ţ���Պ0^��(m㡾m2��j�IZaiA ���X��a Y�~�xJ�q�9��J�E�Q�g���%g���TnoB9A�%����De�_�]s`�╨�`QP�ҍeϝH�������mËv�7�ه��s���٨�&nN�u�~�]��|�!g*!K�lm!�s ��`�u�8�!��Uom]���9orx�tz����2�V-�@-?s�u��ͨ^r�X�Ŏ�N�7��;Th{9����a� T>C�a,5�������nj�<p|�&P������u`�z��B�� ��b>]�;3�4�=�%ʪ�#W���ۮT�r�9j��ʏ����崄H*�	.U�I�1��;5��~�1�(�<�FV8=R�6.��((!hg�$�[�n�?I����'9�M���S�S����%6��d���^i��	� z��4���%`�5+1��1_��9	� �=	�y�r9W�=���.g_�"� XPcd��:R@�!]���m���C�ydm|=R�[��?�m���Շ�Z�5$CUOW��\` �f겻 �fE|sqgS��<#J��ۈ7g�����)ѽ�	��!}9p>rǝ�R=��5|��'��敃^-SRB�)�ׁ����V�-����ޜ�x���}*8rҲ�W�b::�n��+���4�!��*��(À	<�v~c��TtMS%cא�]��|fj�>%�Uyf��VX�\���d:/B_]��	k���v���g*�gry�g脰��*�Ə��P|BZ��]�� ry�ч�r�-��=ؒ/��X�*��Ym�IE�o��혂n:�ǐ8�2Q�!��狊z��Bc�;7�h�9�>�M��׎Ɛ�tg�̛���)=�@���7rz�ųz]|�i%Z�Ϧ6����<�#������gP/��I��lU��sbℬ"/��v��@W�tM]i���*	������$G}9T��:��8e�)��%vQń?������9u� ���{x@"���va�! �o�ٌ�h�OX�H7�l����8�0TF�+�1���:�F��8.Hg��t�:����֮��,=����.O�s�̰o�r~:/C��'l��W�����gN�zٶB�yԳ4&2G(b�7��gP��]��H��&t�r��6��%�c�?��Yi�e�ѡ�jXWa>p�� �1�Q�0E���>�6�j�~�Gs	T�c�>^$k��,�p���^I%�UI���f��\LS��D?���8(N������^�ge���5�xݰ�%)���A;"bp ���y��� '��9��#�˩uu���x]q�p�G�|IH�K�X��S�B�z���V���پ�}�v4�s�v"���Ą%&֮���u-�s���\7!��i��Lw��w����w��5�=Y�C���2���1)w:�_<�Ã�2����p](Ft��J���$E
���j1�4�jS��D�k���"�zMu��Q�����K2�0b�֑�_x��)#�B}�2Fa��HBD!ķ�Ly��Pa@�c�țt,K4"���h�z��r4��KB�Q�Ϭ=S��x���(D�!&E���a!�\�ҷ�jh�/��_4��3�~�!M�W�EL �g������l��U��wUPo*��ˣ5��m���Q�����E|}3�@KNut"3�8�u+��~�=MX� <�̵(�+aԿ�?�]B��u���٢�2\G��,ɽ�h�SYj���|��'����'7��̰��rUgC���Y���"��r�4�C����P?��duS�N�IE��$���}+L+hC5�����B�5��xCv�ZS�8�S��q���汘��w���[۲�<�CQ �L�0ŵ`�>�(~�} ?;���u�m!���xF�9>Y������4$��ԉ���6P?�Y$r��
�(�a��:��$�YI֝��y�h$D�
̂N�6��{W����R��1Qm9��)�r�v[P}��,��5"c-��?�u�� 6/��y䱻��(M�{t�x/T���'U����b�*��1]>#�<�.Eg����L�Yg����N�\=�d
Z{b�й=G�c���|y��Y�J���_&�i�����tx��m�H�CÛ�ah��7��E�`�!XC}��QH�mJHTU�w�Պw��Ȭ�rXE���+����(#��S��FW8庰�G��O�;(!H(/VC�k1��&��a2g�"��~r.��#���r�K��j.ߌ�0o�2�	��v�9A�	��H�B�\�]Ħd^g	�g��k�U�Y��X��G�!DL�7ќaa#�R
��P'oW��1�a�t�6���ٗ�N�Ɍ����BHG��'b�~��=+f�uj��}K0e9���0��:9�����t�i^��>pbw-�c,֑�ux�.�DZ���hG+@����¦xȚTsY0�)]�e�O��G?9�!��b��U=@�\��5~�f+���|Mj2��Q��N|��m�&�a~�-�gi`8�n����<y���������0@�I3o��GM�/�r&�dk�|f�PtG�o��}�:��Mw�K�w��YQ�:B-��<��0-�+h0@�	Ao�N���v����P����f�j��\��ᕭ6فK�Laj�*��J�g�^��
r@Ґ󆵝!)@������Z���nq���Y��4��u�aM����\Uc^fj�),��h�qU=5fF�zp���� �;Iq���ih~W�Qk�Yt�E�����Tt 5@.c�$��O�f�B � ��R��V�Z�i�K7\��<$� 1���QAV�vc�iN��A9���>�������f��U!L��8�э�S2rg
��S͵�*S<���s���$�����x��~�I�BX������}8�7�]C6���_x����0����a�R��dC
H��vod!?��Ւ̫� 푸�A.�����
��f�ʁ�|C��Y��)EV'l��3�W"6Uc�A	Q�H�!UԖ���jXu����
'�-�Dn5"Q���f�z�Z��O,�d��'n5�Sx�<��w�O_C�1f��YT�5J�E��O�q��E����.M+�؉㹧���\��`���SBA7��sh �hbKc�� s���~�"ہ��MJ��֠����P_J�"��oc�nz�a��l��9j;gCϜ=���5_�O�T�;�l}7i�x�q�̪�,���̶p���S$�MFT�����\Vw$T�����\�6�����$�~��;�2f@��hǷ�!��N_���pnm��ҧ�\�W�;��}X�	8Z4���a&I{P5;d*9x�&/=Y������s�j�_n�j���N6�Ĺjk���%�����0>J�K�M�d����
��J�/C������E	��*�ZD����F����lg7
���1$��S�D������&�w���`���
��Ec�/��05�llfC�L��b��:��Z~�?g빫�<ț��O�h"�Aϯ����x
D�B"�����A�MӀ�-���5:�I��� ���G\����i�����n��,���`U�Oq��DMx7��<�c�>�w��yq�{�hr#��!�CI���f���̰
{[k�W�N�e8��8�̠���NaӢ��e
���0��NpEV�"�@[�Y�,����G3d)ҬH��������o9ߜ��{��n�ر���J���ێ/�v�E�6�= w^���:��S�(����8���8�D���ȣ��<f�:K{>	�����;��Krx;�?0 �`T�)�QU��ġ☫_��*3˙���������8�r��LT���w���=��ɤ�}!����� NA,6�z��J��ctt��������h�30%{������A#��"鳋G@��?��	�u8.[^؀i#�r�-�f/��%Q�eWR�B��q4��MH��?��SN�C�2g���m���\��FoK�m��<��uׯ���JZ����.݅�
��Z	$	�ň��cr�p����o�O���bP*�;��C�S��7�<�J�p�;s�i=g '��F�Q�b��ٌ�|?���%#%J46i!y��ʻN�t�ZfڐH����ؐ
uk�Z�B�&/foغD�!�:f=�9np#�?���ϲA�bS�~I�^-xC�*ڑc�D5oP�C��2*�^D?b<��v]�{�L��y�ژ+d�R��\�>�xǂ��b�E��fF���h|I�wEԂ)��w[��A=n1��.�T��u�hJ��ԣJ��@��ń縉���(� �ԭ;q)Z�`�n%��yRkx��� �����ú�`�
�Oa\u�A����	mmF�6��՞�'�!��@\@Mi�:0�!���U���t<۱�@�,��֑)uD��=�:�Cq��<s����F��Eb[�7�G��!y���]�*�Ț�&��i-�kW))�Fd�`�(�7Q�V<㤷��mo�Ӭ�݇ؖ��>��Ӵ���k-/(��
�b@@z�&�L2�|�ЏHگT������-�
�_�M:;c3�M�-��S�r@lǗ%i]��g׍d�I�C~P:���7B��!�gg<	�݃����������GVhf��w>���1[0m�%+��������y�*I��mW͡x7�[s/�{P�i0�sV����͈[�$�C$�m#0[N��cC4C�?�Z�?%>bF �i�#*����]�+kً�cd�4`M*j>I��^!)KΙ�*�r���H01�nҊѹ��_��/8� �;�Uod6-p���V�{1���ԡ(�`c�'qY/�K���݂j�;u�vt@t�G����p��������$n�P��i�zJV��?��e�ha��2JOn���\Γ���������K�禝Ƹ�Mn��=�?���8s6� "@ij#B�6��;7�T
gc��(g�x(N��\��ÑV⅔ w/t������-�2�y�*�_z/O�+xj����l�Ut�������~�=�8���s�����A�TS1�_����U�~d�"qH�+n�_�)7ϒ�][;�Ff1��>��O7�;f��t	�s�'�.F#��Sf(�:�·@��9{�A��q�+�:��NY��V�KѨKg���B� �Q�{9�����Ő���&˰�O�B�yH���"��[W�<0��t�k�އ���,�f�b���]p��=����e25
�pݞ�����^3������uNۦ��]a|�-X�iK�n�˒�8����+M��0N�G��N�sY��9*����L�F7��O\�uuN���i~�ja}�,pby:�;����`ē�u�.C��!Ez󒟼+t�X0{X��t[s�ß�yy�h-mM3#S�{�>0����O������(�)�l���9/"��&Ғ2���J�O�$��1�0ҭ�2����������FZ�ƨ��gy�M ���2�@e�n!<����4��(�5��w}�lĶb�q#!)�*��f%��#[sO��k(������X�L�ؐW̿�|��������o��hS���U����d8*�&�[��r<��V��'{`,̆�;@����I�[���춤��`i�%XΙC_�s�I�q	E�:4NA���c�
ٺ�gA3#���
X[c��:ԭ[�	W�l���˓��"����a�r���m?��7�A����E,!��!Gp�+@�'�����C�������vʖ�3�k'���� ;��#)��v���{�����#�hة��-�6#4��pK�U�oS�e������8��s�/)ֶʤ�7D8� �NO|u+zrт��S�6�ȑ�>�XsPq(?���m�������IK�#����k��>߇�Π3]�v5��w�7��s�P��䧡�kd�7�v�;aQ&M����Չ���Yǉu�����q*�]b?��W~;�����3�t�ˏ@}Y%��V'37�ӟ�&�5d	\��%?���8 Pb��[5�U&�vε!���ڵ�����C��MX�]�q���e���髤��dA廝:��DI��s�+_�,	b�
YH'bEZv	7�4����.�͆ϩ�~g�	De��i=��y�j�����kr�͍���b��W^_��|U���X	'�֢ ���_�t�Ɲs��#�&�˙�j�q3�{]q�[b�r�ϱZ�,i6����#h[e�oΛ���*�<S �,AH��,G�[����:S^�j���.澼�`����7V�j������cX�)�RG�`���SX2�6��&�8}�Aۃ�T�QA�&�
;E}nnD�n��v_������0a&��47��C�U��kX'o�d���b����΃�Aĭޱ��8����=�B��UQz�?��R���8�)�z���ko������у��jʳ�XlH����������tb�vr+�8��"�yޏ�3���D�-
�ĐƑC ��������EW��	���o��K�i���M�TI֖5`i�2��_&*�?ݴ�����͑�O�A��+��].̶����`=�Ha}~MI�,rhsK;��K��R��ihC�o��A�
 ꮴ��c�}]��.@�,=�-h���j��������4W�Z�mIqu���b������Q|^�KB��n]%�S�S�hRO�L�_��f����w��`w�? V�:�c>[oouJ�:��l�o]�Y3
w�z�m���24z�OQ)rz�5�Z�<m'=���򟏄K��IQU&�-��Jcb��i�i�a�4�`�sա��2�bk�rq�� �j���F����:�@���<z�5rX�`!�E�,!��d�-��)�����`}"��5�@�Eݑ9���q�m�*t7���
/�e���J��W�(L�Z0B���g�2��r��-������
Dϛ��� {��M��8�r�u�p�¤'{z����!i�zsU>�^�䷬S3�l�� ���짭������,��^�2����p^&��c.��
}"���	3ɠ�	k^#G|%!;��ep��"�͑���
�û�+�7��5�H�"D�q�9�[��<��G�#��&��z�����-Ep"�����'�N����:�R@8��v�S��^�'����B��YF�ey��^u��������t#؜�_������v�*/;�a=�y�$���+ԗ�� ��#�7�9��I��<���ak����� Y�����ysopwP#Roe{p� S>)#ti჻�Kh_�ؖLO�����zÍ�X�"U��4��E媽�k\��� �����/	sK+=4G�jF�������l�=,�Cd6D��O���"ЫO�Q��%H��jj����eW����QL��]
��V¨MpQ�7\�ﲿ-��]�e���%��Tf<��?
�a�z���~u��"tN�����#~l�g���g
��X��_qb`��������P��Pysaf�|��?�P(���0���p],)ƐE
�T���SQ{������5�G0s�cq@��Ҿ$���uM�lD��,�"�5����	�攞 ��:o��ֳ�=�%�;[g�P5�獺�WOW-�b����V��ZQN;G1��D�Zc�!</�'�Uy�)�W�(>�k�����&�%��
�ͨ�uw?b�</$�1]����h٭[�}����4����&|��%�bJ���7�h�t�<���XѸe��Ym���&��Ǝ���`5�7��[=�r�����s�C�k�9�ݒɛ�����4����%8�T�-���[�����/Ze�C_�)%�̱O�o騭�)�l���Eu��e���3��C��P3��+}{��%W�������&\�n���)���Q�~�d9�_Zs�YO(y�E@N>��w�����!Ӳ�9	�*) ��ciýG�����6�+�2���hO��Դ�Wl���SZ��[XS���e;[�[�#yc5��J{$�L���� �[���:�\Y��߱�)���̟�6کy}ysʺ{���x�,�Hhy�e�p.;>�J XV$
rwغ�&��3}�Q�+"�C�� a��*q�}�O�2������^�	w����ئX�������G}�b?�#TM�H�N�i1����n�I�RU��D��o���HC�%��C{�
�")�g��Dz'rTs&��@o�)��Q��0Q�X+N:���(zߧ��8�=jɬ��V��%}z�[�1��g�?Q����%�q@�#;M�L��$�B���^�5�ʙIT�l����7F�F�Y��*ds��sC��e	 n��L�����rkE�� .�1G1���g��`����1�Z[`���S�b��y��Yu��d ��N�ه�le��vZ��t�]�۠v'Ȥ��U�4�{zsv#|�Z�����|��Ŕqc�Z䖵�w�[���h��a���Y�V���G�xD�I��X�#_�v�&kL�y�F��օ"���'�@���g�L�b��z�`�X�'%J�OE�(�nt�}u��!VC��������q^�y�ӆ-�l]>j+M����A�Ɨ�,��`�=V���1�3�*�4С��\4���u�НZ�&��(��f\n��)1��
ġhb��-2�&��!���(<6-�D��y�-��h�-K�2�&�v�F�_7�@0���UK"��_��U�	��߼��ރ��az��H�d��w���#^�!iG�K -����cR/9?��u�L��6٪�7]��y���!�ԬA��R���g��\�T��(��.���?vo~����	�@H_���k[�鱱�yi��M��u^�R:�Kt��������,%a���qaoGb��'�Y ��sxy�6TOd'y���iR�����@�7�Z�K���P�����*-Կی���ǬOt~dG����DP���ᔩ�^��AB�7�H]�'.5iHȫ�8����U�*j�1l=F8]��c.����=�����,���E�g;;yYsC�������\�v�|��n?��=s������Cց,�����W�X���^�TV�/��A[�s���)BX���S�]Ta��(e3>�U�&2�,D�̈́�0F��/؆j
�@�R�}�6M�]M�9�1/^m���EdT7��d�h#,�֠d?�R�@i�M˿L.��Ɵ�v�/�+Lqiʳ�^�S�l�+��Ś������L���2uW��a8���*���H�n�uBe��j����g�I�����i� ����{V�F/^��:t�nS��.���u���T^lڛH n���{� L����;Y�a��uo���cL	E��V�C�*&��d�c��KȗR.Ʀ�#]��y_"?��`��`eF���Vb�=*�	Ɍ!�}�%2qZ�[��p�o��^^�ɽ�J'f�� �0^�U����[需cڷ�)�Ҩ,iS{���|a��9|�*�DE1������;�,-r��hʽ���~�^Pl�Z�2P�5���P�-���h���Q�(OP kȵ_�٢�*GCg�)�����xç]�0u*ǁ�$E���yՐE�*��t�Ǩ�S-�~�`K�BE��*�Sd��OE�M�IP�rV�jVo�t1���e�Y<أ����{ʹj�gr~���̱JQ�8a�*��������v����� �ޛ7W"�>F:�W��g �L+�R�]��{Z�c�T�ھ����gʨ��i5�
�G	���v�F46UZ����P�� ��Y��1M�e�;|�V����)����k���X��:Ǚ���G���r�����8ˋ�9?���q^?C^3�Ru�B7#�?��5Û(i5*&^�İ�G��_�/��K>���$4�+��L-��㴫��O��!�ץ�0x�Tץ��>^օ`��Y=���yU�ZJ[� >
9KҀ,k�`�9ɶ�z�˙�4rL�ZjBxڢD��>O��'�II:<89Ъz#�~`W`���{L�r�v��MN5��dxa�ܫJI%��"!�N��(��'���I�^��U�����?�L}��&i���ѷ2�����I�K�2�Lnƻ9�%p��a�?��m��=\�5ųǿu:�;4�c����ȅ[�ǔ�s*)�t�\�j �J�!fά�k ��o�+CmoN�����Y�)���-.E��2��p��>T��_!����-|`�+����c.⵷�-z��W�eސ�ia������v,����2�%�0��޺E���Hт���ٿ�=Sz�����J{�.�d$	V,��#6"*8u���D;�!�����5�t��Җ:o�=���~���ǁ.��[�ڸ�}1�ߕ6b��J�x~=_KX�����~���]��Pٻ��G��zt�o�k_��Yqx���|T��i3�B�&�`�;D�L)�1Wѓ�.2i���&� }6�h���q�R��R"C��	d���f��g��Dr�Q n��Q���(��gi_-!�M<Rt�ή�5��H���WU��%E��Us?\��t��ɿjk��؏�o"���[ͤ I޴�?�'����T@�+�ݛ%���z��?-G�%���ic�|�J��F�7�!t�Su�7�<7LJ������39�2���IJ��#�[�VF�|���!4 �Ꭴ�&�%�_�Q���
��?�C�?�5���5"v��_z��� ^��(R�x��a�8���V6���������ى��M@.�񼢂�v�C�h��8R����1�3W:1gI�^ ��}�������wb!�'ŶRL�,s�dG�mb��C=�(լ�|���쨯j�
{@��,�o<��L5��+�Y�o��O��,E����r�ɍ�wy��ɑnP��#j�g\Ӽ3�{�.�߽6^��E(Q������1r�\���wewK?È�����F�i�-aKk�55��<�Jt얔��k�$^�Z�-%�]��Eg?*���A����b�=�َ�&~S�1 �i�<~B^�z����Öt�ES�#jfc�ܙd�x���c:?c���w�,�M����zǫ0�����	�L�����{j��H�P�˶��|l7v��{ژ�'/k�p�[P
tU8\d{��]���j�sj!�\�oc�O�����J��"&��h�P����Ǳ��Q�q�S|�,�Z��ʚm�	��r��V˓Z�+!7�`����ȡ�cS
P�h�Ľ���2OM"� y$�C�i[����@��ȵ�R��M��i-�Z���N8�t������Q- /���]y����s	@�!`+��GV;���[%�����S� �����8�Rڜ�kP��si;	�a�.��0��6rZ��{����&i#���
)��P��
�=�:��D�l���c�����r�tR̳��Կ���r���+�M�+��hW�O6՜�FvX+����v�b+`C�t4��5�����;.򎠠��k�z�#� ���W�#�1?����A0utӣ��ȍ�WLJ��lː�U)/��N�m%���`h�5�P��^�R?���sYFv6�J�2���h V?�Q��,��Ԃ�v�!�9)O��x��TB�	�'1��Rtd'$����q��^�4��(>��܍�tݮGx�^M�Q:a����8���ʔ�JB"�V�3ς�����/�[��CH	��A�=��rя\�)�(u��2�J�9��O�z���bb�9q=�8��Q��i�	=��K�Q������>h���I���ʰ���f��/��{�-yF�~s��[���<��9?Z��֠l	!	 �[�R=<�ƴ�©�
�Wj�t��<4d�*G㪫�4�	�e.0�(�+��]t�ޗ�����&��VŽ#���.���@'m���u'km����璼�,�8^f�c�bjR����Ǜe{�O#_��|��CG9cdJ7��@]@�$����.׻�.�,�U�=��;�pδ���ߛ�"�kT����h�<�qS"ʰ�Nv�zy$o�T�_�4�&��C��W�i���ЫK��G�;�~�oM���K���{Hk��!P�:3��V��Y�S�x8o���S^���<ZB�̠|H��<x��_y��d'`��K���Nd���P!2�n��"~.mp?t?�#�$K�¬�^ɮ{w�j+�$g����8��K�8_A(�W�)vK�|�b.C������ G�2����VJ�-���Q��8�	P��7%���#a�A7��i˱4G`
-�O���2qÐ�$̊�)i�{��u�i�f�P���&Y�g��#�x�NR=��tk�'�x��+a�y����Y����*��+Ʀ��J�0^s��x3��t�	���8|���hǽi��=K[}�S����C<��05e���0PjA��K���kS����6�n�:�CwP�iO��xIN2l�+-���8�����X7X�@��V99�Zμ���8[�;<؋�����H��,�8`^�bW�����I>��1���ة�p��ꔫ�j����C\�	�ց�=��{�нÙ�D;�sNp��|�S~���lrN;N a�����ۆ��쓜��ێp&���܉Gk�T���;�[ˌ���5}�7i�3XM�87>G �H<�Pd�1�}l�H�e�EM;����:�B�Da.�&U4F��!�g��C�Z[�N9�h��i
[v7����@���=�<d��[Yi�q������%`�ǒ�jLçGFN!��$�^��\��q?�C�M�*l8�"3k�OAp���YlAU���F�R�3￠��� 14�e����n�(exqM�VT`s��h@ML�Ġ��Ө��<���p��F�5k:����=��X��F�9{tl�J}�bŚ�?Y��j�$�ڧ%�l�A���8���{[�]I7�d�"09�����vm��]�E����9�q�Z*G��k���:����sUo-��7����Aj�]�V�C���.�dŉC*ɖ��E��1��ǳ��'n~ޛ��G��43�1~�B NdZJ���)����P������-��x(
v�����W�f�_�?k���;�?|�+l`��*(3��8W��k����g�������&����&~����V�9�H���*����F͙(`#��۽i��n؈�R�Ӽ��Pm~�{g>�AG�S�]u/M�h��(��O�8��l��0�SRR���)�<Yr,�Ph#B��������H�b�l%Zz<���~���Rw�t�����ʴ�joLp���86�V��у��$9a2D�j��ȎY�6I�ި.��9u 5�c@�k�s*�8iV�1@�!I� Y�8��SN�}yHk5�A0���B�r`�Ϋpdm��?��>�?�D�Fg���f��(pS�Щ�M�3>��KjUi@m(����e��XD�}��ϝȪ"g�	����YΏ*S�����0:rHå��}QP���:(�k��A:��:2��}F������z�<��V���O��OӤO���lwx�CJWP�]'$���������ڠ���X*/O�2Z��{M ��"_�?�7� #���VA��e� 

�a��s���n8�I�#^�}��@ w�`��̀}�|���c#Z|��-�����IRo=�����H�(�0�O�����V��<����^�&�$��
O�">*g6��T&���p�ע|�:x���L�ݭ=�JR��~;�Blަ^��)׺V@��j�F	�G��zp�Q4'j"w^���U^��s��`c���� �E�=]$��������oԔ�cȚCї6t����|���q�����K7�@��,����Mv�����Z���At��m�@o�TJ��G��b�2ٝ��r���f����>�k1��jn�
�cȎh�g��0GEu���J�d.�i=�G�z~�Q1�Wq�L�)����.�*�k}����x�l�N���R�X �w�f�>�hh�z7��A�G��ӿ0�u܇+T�~]%�#n��xE�wGZ�?R��q��ߚd�e\�jv���_�(�-d�ͅ��7���D��{b�aH�]�ՓqT��+G�(�d�W��9x� ���S^GQ�Q�D��K XoP�&b0W���C��6�]��D>�t=�D��O�� ~�N����B�?ܤ��(�����V�
e�T�K�x��QUǨ��](ۙ�����T602i�:�8�{����C��Q/���0l�T qZBp-��$Xj�N]C5"$%��H(,J�=��_$�p��^ϥ�@���U
'��Μc-�C�E�W���9''���.+�k��T�jc���-#�		�QCl����mW�gB	�����>�ݕ��7^��z�p�Pp�s�޻V�B�;y�I��RFe-I���b�h|�ݨ7-�g�&���R�_�Y^���C.`,�(�2�۱r�dgʔO�?�t��>`SG�	{�ϑ�j�TG+��D8��&��y��>�Өd&-~�<�o<ġ�<RAF�X�DML I����.���hC�	�Lp-'�=Y�s\�e�5v��y�2t��I,���[�kō{��߸�({%�0|��JGg�e�����K�j�h끵�"o�O�]�4&!�C�b�M�qCҔ��$`�|��x�����Č�C�h�o��7����3�o?^pJ
�����ǖ��$��̼�>tc�L���e�	��i��R���s6]嵄ؼ^����i��QM!�o𣆚^��N��j
�����`c��Q�IU?�3G쌜B&�w}�=�����^w�8�*v�����&3����N�y)�3�w�L!XI���^��ܷ>g��$��{���8�9����ܤ^7�twҍ�"�J������m��V�z�[�:4:���qL�T�o��3bH!)J��G���,�� �A��/�+���(b{�'C����.��[4]�0*�<�$�'0�����/y��+�m��d4�f�9�B���N�/���8BMd���.c�V3'��X���%�WL�3�W	r
�ߎ����L���DH;SY�-�7�/O@g��p��:�[21�cG���vS�en`�v��"@�uB I����&���� )2�φ[�!}m��}����!���,F-X�c�է�� |�$L�aǦ�%�ݶ$?��&�q�����|��j��{�ڐ`�9g�d����N-��{sUQٴs�;zՏh�w��s�vT���#�)���uN���/
Ըȃ�b���~_w��<�F#2��8>�|L�L�ETP-��l��0�0[�����Ռo�k]��[I�5磉F]cz0(���f���N��5L�H{U\i�Ь�f�ߖ� �a�(�G��"WPf0�Z;˖|��,dY5ܮ%�A0:1��c��,���=��h�W��B����!{$Q�3���N��U�`��y� �T7:RF~J����� �z�@j�D����K`%�,�ؙ[������\�ɶs�S�ݪB�Ï.���I��G4���$}ñP{䃅r����[R`i���_A8.KL)R�����O����J�"��
J�8H�� 5\��Q ��S2��4��E݋:��i�NS��=���6䅤m4�>.jvr��%�Zj�AZ����x� /ಟ�a���vZI}��QpF9� *��ktP���u�Y"1��&�E?����i��b7q����R�T��n#��_=�l�9C4<=�7Ch���_�x�+��b��~�Āە0�L������כ3�>*��#%�^�$��p_<�(uY��h�w�R����X���(U�ʯ��\	��L<����NJ
}
����:�˫)��Br�Y�g+�u�Q�\COf)(�6Mؕ5��H����̍]�
�Et����\s��zp8AQ(N&�^蓞���n"�eR��(B	J$���XB��,3��OP��@��}TZ���O�3,`��˜�\�9�z�L8D7u��s`��$�Bu���t�I	�T�ey��oHP{�ϰ�'IJ�z/�ݫ� 1GcH%gsp��-�G����뙓�2�#����U��D6l��ƍ%�
�4�<��i_t`|�C�z]\�T>o5�Q�-)r�G�l0
�o?ڴ����G��^����M���$�(0�oacBAϣ���]�<0Ż�D?4�4��(t��ƽi�_��>�cM��5>(j�s�<��(�TQ*�����߫B(3�lI�g(f�W����	X�t�+���Y�7VA�$Ƌ�6��i�Q�3�9�q��d.[��C���+dcJȇ��S}4e�Yb��e������	k�P~��VnL������O�����[�y����������Wk�U�ء�Ԃ�3���X ���3([3S�9@=�ײ��m�"��� �غ����jxs�ԣu亮U���S��gza�������i�W$2n��K�,�+.��8����% DGZ�ͫ�APp���zJ�S���S������';��L�_��N_�����,
�Be�(�X�>$&3�஗��=�B�U,|"��,C���kG?�m�Ԛ1���ll�6�Y��������Jl�1�Ř �B~~)�7�?K��sIh�S裧S��;�&�<�zx"}{�ԓ�ޥ.�CpnAֽ�E�Q����6��ݖ�d�C5����h����M�0���[��a%	㥕1�:ș8i��k6�� �i���������@�:}�c�%�HU]�a�o�5�Ơ��o�$���� ��5w�3�)�����b��q�9��fE}>e]"qh)�?����]�Y�I���
l˛�XCy��Q���	6�o*J��h����%�b���6p}:�F݃˘�Jﶉ��p1�	�p\gbW���z}�<��ȓ^���u�Ecq6:S$E���x�k�8d�V��ldaU~��
�ɛ�2�e��V/5) m��j���9ץ8KNU7��I,_�W�p3u��ר������~�����&�I;7��\��&��E����p��W�j��R�)F�F��#�"��甅D.ǲ�mNq�'������j���sJ�ޚ�nR����S�JAS�v�V=�Dtȹ�4�>(&������%�����y�L���!�=%�le_�Q|#�nm� �&��u�S*V�H�-;@NG�q�)�����;�	E��AVQw�m��Cy��;��� FV�	�r��֋�C"}%3yk�+w)ꙉ.��,��Iw&),�<p��������f�#��ߛ��.0��=�aR�� 	7�Ge��oh�ׄ&�;g5ƒ����������Q��*�4�I�U�P�=o�h��`"���}�L��*!�OU}�Z;�.��VVS
�3����^���r�Cs�����"Ʒ���G~ވ�$N�[H����](N�NK�|k���)��q���֯��H�z��O�7�䟰-�D�^���8/u�A>P��߄�<JZKI���K�F�Sj�󬫬���V�&_�<Yx�u/0��r�;;���Bs���윛�a��ff㓼9����r;҇�`i��t��fȊ�c���I�?6Q��Wqe��5_EQJGȚtA|�}�7ֈcq�"P<Ra�Lᨳ!B�r�TK|Ds	��h���%.���h�1�'���6���G�����F�/�Q�G�jQ�:2,8_w\�G�|�pzD�R*��x�h�@o
Z�:(#���c2qm��r�8]t�'�hI�@16?j9��+�N��8&�-ǳ:�K�ۄ��|i�!RO��d}7t�r��XJ��0y�a��P@K��P� i�=��������G����yH4r'�B�������?n�4{���v�s���:�z��L_�����s��w46Y&����7"��� 
h=^Ѽ����`�z�C�_����<�ܡ���oW��n�,�@M�W�h�L&��`��/a�q���?�z|g �wJm�@MYԩ{�����eq(p�%���3�����K�We	Su�%a���i�������-u.]CӤ�!���XF4�Zy��i��?{��,o�9�������F�c��,�x&Z���56��<J��x�E����T|Ň{�un7b32
;ryE2��{�@jZ6�%m�:��"&�2!`�0��cr��Is�J���l����vd*L�`4����2���w<Qc`�2l���B	$�3�!1��a��h��#��v��鳒��lͼt� �󊫗Yt���j���b�M(W��#0'X���娯�~��!.YÉnx+�� �3�{�)�n��NZi\1u
���n?��;؟Z��ka����_�ʀl�����oer�?s�F ����4��%��Ĥ<k�t/6G"�`�g/o���*���m)� 
�şF�oH��v�����W��J �g_��Ʋ��Da�CH��/˶�)E_鶆R;E���*��:C���X<a8��pI�Uז���x)���"t�S_���(<~=1?�X�b���"M��L`�)�ݵ���|l����M,�`t��X>�j���pKjGN^������ʄfmr����a�Z�nt�Lm��,��෗�5����m�O���<���pBꯈ�Y�*��7��6�}	P�� ���g��_9K�t��z�Հ܄dLxs��ys<Ψ�c$����&';J*8��ƍ6��ZT����kШ�c�khS؈"��B�� ��n��g��u#P&
�f-����I����:�G��Y��P2����ӊW]vt/R��WLn�=�X�MPY��m�N�G�Ƃ���J��[�H��!��h�~��I޹s�Qc�]Ԃ+�yW���W:�-��Zʱ}E��C��Q��Q^#Z�$ ������� NШf�T4X�M�c��އ�X:4�ʝ��us� ���Ǫ��,�ob��b*���s�5k9y�v?=g��|*k��p���ZI�Wt���@��ՇK�+�G�D��{>Cӯ���w�Ω�$8����n��!��{�� �Qe)N�o�Bc|�s=ʷ��B/+4�	�s3˾}P�WY��љL�v���zٚO}VwHG��V_ֆ,lz=��:I�C��G)1�Ū�To"�����P~熗�{ڱ���;�U���*�_̊3���p��GPS~S-#�� X̋�cu��*�-��D����T5���nY)rX
�>G��s���^zo�aD�o�
�RW��,F;�#`v ?�� ��9Z&�d|��ߡ'�W���*�J�����C~��&�k����DS��C&����o9P�2�p"6~�*���%�a�g�� �g@��c݄��fO<��LΕc�؜�����E]�,���u��jlN��	�7��w�q�j�Z�0z?nV:uJ�sV�5�a? !v��C
�8�GC��T�ft�jws\Y	���m�sň',Gp^�g�/[�1��UL9�S�ᮉ�e��c3At,A��?��t��w�vf���g�
��x_���3�ýMq�t,|��0���le�L��"?�n��nY~�x)f�!oA�Ի��ns��%��8������P�b��������������/�yIe����.�U�����>�[��?��ߪ��9Ha�4�ֻ��{e���(�b�Un�Hĥ�8I,a�^��!f�=7����̧flSF�P�9p՗Q���#��R)|�%gA�R?I��O e���!����c�t�7�LkmR�*"G8���Q^'����}
��6��CҺ?��eO���k�����
t��H��B�>�L�PM���� �hAXT�<��#I�$�m�Ɂ}K�XC��H��`�8�,��N�#"������+��w�uO�O =�7�#�����;��[�͸ �"��z�1K������;o�e�RG�k�94@��Ԅȥ�{��ߊ�����J�#��b�zG�rUGv�+�1��rQ9 ��.����{s�W�{Nm�k���N���#��=Zu�%�v�%)~�+���>ݨ��<g�4wa���S��L&���2�z��5͋���Y�D�:�꓅��V�ρ����sDu�}?ק
g<���ρÜ�dq�C�
��p)����p����\Ij�z���\+��yLfߚ�IK�|U��.˿�P�[t�#n�8cT�z��%��3���f�FP��\��c�z�&��oG�a�@�-��f��,��V��(�R'tt�F����F�hq_N����c�s8�_�����U񉱂u�~��Np3�l��'�oy�}��|t�e�4=	��k���K*�����C��X�6^&�W�T�Owt�0�2di�n!'r��&%Խ�X�9�����PF}W���H�/K�	��U�7�Ed�hT��?�sĄ�7��0��
��؟tw�pE[ӥ�~�g��s#D��pc��ܜ����k?d����B3w��r^]�Ļ��*�\;�˝&��1(�Y�E�hm�Ƚ;�zl�8x��$�9�
�#��t`��@ݦip{)�J �2.�>��(=��?d��/���>#���0�׭�OBd�L�C�;���oQ�'}"�@��\�wȇ���
��e�	 U���~��0����`�aY�oa4T@�A��1�'����o��oQ��rLx���@��%��4}��sS��r���H��7�$�<��7�}��^y(�i�2S�\=^�U%�����LlX�_��'�C�-~ψ2~ՙ�*�F�	�O�������7�K��0�\啭�D]���6%������
���H��0|�ܩ�1���������%��R�I㖲���{X'���
j��Y�=8А�WQg�A�.�hi��󌉃}�e2�;�!��p]b��@z�ݖe��!�u9�@սÝ}���$�_fn\�g��a�y�kR�\�fh�����GU�V��D�$EQ����t���g ���U�sU�RQ�;�5;��*�Ŝ'�PF�$V���{v�s����5D�n�^��wx�QoŌM)s�V���RŮ���,��0�H�k1��PM୆Y���v@�B���G|q�\{�OE$ɒk���m�~ٔ���T[vPѹ��N��|�P4%MY�>7�+q�;d��Lʧɻ)���]����<T�M��O�K��9���ۜ(=�{�����������͘m��$$��glhDa�Jy[����ps�-% }���&���ҹ�K�x_b����$�*�-��)��vP�o�O�G��/N��K!X8�Q�6�H���5-�_��!�u�u�2"�;[����>.�$xa���GF�Ax�;���صT�y�0:��ū�ߴ��ލ�y�ODO�+w���S�V�Yw��9��*�K3Ґe���tf��d߹$i�[@�g���#j�o{Z��R�"��@�{1>QA�M�"qI��̰X�!JS�̳��C!��n��`T;�,9)���~�W���߾��Z����Z�c"QnL�j=�e����P?0�pf1B[���,����y'����d����U�l���f��������z�sĆ���\��qc�oE�PN�A�j����w�"�������SS+`��ž_��h�ڍ��1N��V��Ɯ���NTb�3��p����2p��������� �iJH�B�V6W�����q3����쪓�降�?�=��uN��3��?�) Y�����b�����#:5� ���b709��0���"���s�^���n
�;1Øն(a-���q�I�Ɋ�v�y��ի�Ʌ�52�s��-Χj#��J�>RYI9L�a2"sT%D��ޞ-?7�%���f��bxR������;񱽀N�"d���["�N�gf�������z�b�yF	���M'^C*��W�.���(�\��Ź�J��5_5Wܟl��=��0<.r���^{�+e_���)������p]_I����@q+eڹ��t,X�n�O���%.of�gf���(�@�Ғ�b���.CV�a���O��%������8�Cl���sh�$�̓DV��&-�}��I$��<�s3�3�*a��8�*-kцw7��A��!�xڑ��ئW��V���<�/�l`I.���5�d�N�TWŠ�cB�,s��y�VPF[���z;�=c��a�(���.v_�<�|�m�u�d��b��#��^oZ^D#	�_2m��rp��t/����׈�wY�(+5V�,�r� q��ڝd H[�N����qI�k]����7r^f��?�ig�y�΁��|i��y��o!O��!>8>}������&�-l�i��E_2?ȩ2�ɭ���h��״�F�V:�AӮ4���ځVǩ�՛K$���x��V։#�t�t�vF&�<4T��vL4�d8�^t��qh��WR��e�ol���S�vc�3�8K�Y�����L~��8��k�<J#`T���5O�Eb�ƪ?��`����#v�;������/D�m|gb�訁� �ӷ�J��������L�9�dogwT,y��1x�ҫ߱���� �oKGL<:Y7�ڇ��(�N��;��l�͌l7��	w� _�5&D�!@O��9'�1�Έk;��w���?>��e,$3�G(�@���.�߲4��k�j�&zc������i��m�u� k���-2��=y��Tv����S���Y�&�3�"�Z/*H���)n�U�ľ{�|�c܀(JH�k�?C�{Ȇ�\�P"�p3��P����PUk�\���-¦��n1�*a��{[�م�nP������)����N���<̻$��&��w8}n�7c���D������J����JS�|�CV[�=d����).B/�X��S`l��-xi�	�U>Ɇ(X�m��6ETJ*�5�bx��-8�Ssۛ���>e��^{;��Ħ��-9��r39��	ӏr	�����H�)I�N��ġ� ,�ŃAB��y�O�s|w�<LZ?��������",����9����c�/��rc
�s�~�wB�/$�F��x� ���	O?�c�:MNg�8�:�AZ��Z�ĮD_wUD;ײ �=U�ҧW�
��!c��`�&�N���4�(�s��s�����:�}���2�-����̪�}�=��ȧ.ܥ�o:@ڤV�̘�����p�km�o���mb+��aY�i~�E�J�� ��KD�1�2�=Y\ڞ�	q������dR�DY�20-���j���N�xoߏ�S�'���g�⟵��$��}�������r7lW7"�N6�OJ�[�-�Sw3֥�/?�-�Sqh��qb�/U48�(�ߊ\-��Rt͗���?K��\/��(��d�0R���z�N�R%��B2�p}��.�߈�����K����?�1����/�4#�O�g���1^+U8/�KM�]���׌�2']E?ALm�"���᚝�T��<Ln?&�2��$�.�
�T&��Y��v��Q���/�^��G���~�qAh �� �/�	�|���;�7�J��3�\?C��Gp�W�ϋ��#��Xz��o1Q��]u�M#84��MP��TtZWpѭ£#d�i�)T�(͇�/�s�ɘMs�TT_X�Ȍ]
��>��R2^������'�`t����ResW+l0�	؉*xŗ?��{��Y��o����R�r�%+/Rl	��#I̳�B�(S^6��+�����<r�u.�(o�pJ�#橪B�g,��ܖ�+��$�.(5��Ǔ���S:xG���f����h��ES��>u�XQ���]�����-ǀd�f��@����H��T!�/2�pX�v+=�K6�n!em���q�[�,�(�9�J��ff��C7������s��I��{�+�1���U?�
��I��"��F��Q:� ��٧9��{Xҡ�D��t&����u�u/ aU���W����.��E��Q��N��;Oj ����$G��{�����@֛J���^�{J]�լ9�q9_ΘEmy^%��b�CP(�̦u�i�1��&�h+_�讦fʋGp��⭃��I&$du�C>��`9�8���?�qB���MQ���W�6��켮�|��O%&I��}m݀�Ĺ5Z/��I�|���q��@Ӽ�<.]���Ȋ��߂Xy|�G`�#���(�#���&D��P�YR�&�^��ynh>D=��>�=`����s�>��ž�6�מ��"D���y���r�jEg��8s�����X��Y��l!�I����*7YZ�0���w��@���i��.S�O��$8{̭/~4#���x��x����:�w(���Td�z���L��i��-��@1O�[�0��IL�c���\U<F�}X�-�;�$�~	(t�mP����up|����W�"���+�=ڬ�wl턿=mІ�(t���42�ڬ
p%�d�Òj*�oS�5�^{i���0-��e�j��5W/�����ͷj�ܭ�o$�vF.�C��i��#�BJL(�l�����D�ö�����9�N��9 �l:��G��9ş)���z�$�'���+��Y'\���n�`�S�1xԥ���,BU��ZWQn��Ma��wT�h3$���J��bO�3��oİ�jy<j��-j��5}Ϲ+�_��g~h�wN*�8C��Q�VQ�d��1�1<v~k3"�YZc�K�mn��/˴���4��4O��(�����Ӵ�^�8�d�h�7s�y��^<:���M�'���C/n@s=�J���W���ܯO�:�; �ݑ�^z��`��%`B�s��X��� ���r�,\#��YJ0Q;YQ6���h��㥑��s#\"N�w����v8��ჹ��1M��H������ǌ�v/�9b���+�D��pރ�:�2��Nk��q󯑪.
�O��f��ᖊ�kr�*:6ۛ�����~�^`X�D���(\j&My�
�ώg0�m5�˗���x`�)_)n=����wB0�P�D٣� �:D�f�Y��X�3� �T�[Dך0ؔ���jr��&J�p��a�IDǫ��cO��u���̑E����|�G��t'� y����g
}Mu��ީ �!�9Uf\L�*�w�ˠ0D��b`.X�HY�:�9R|�L(��cн�\>]!�F�bj�ME'��Z��Z�K�A�CyLP���#��,��<�e ��<Oi�	��i���uQ����� �&�gi�ܭ�K�}dLn��d�!A�I�̖�Y�3tp(O�n�>��sb�C�<���>&\F����Nu�(Az)�߲��b�M�qoY}��~�%��螻8�g1���'72�{�'�85�X�(�Qm)`��[:�.��%��w�[t�ᖊ����uY
z�͵�i������Gy�U�K]�GV�W�|�n�/�=u�\ T�XIn̈́>��,�ߊ�;|�:�)~�	�_��nh���F4���)�5�K!�?l|���J$U�z�tK�#���T�#�{dJ=&��w�EW������<���� ����KMʢ�όZ��f;8�	[�&�Hwp��Ș�gG�F>Ca����0z/�&�?�f��1Y�U���J+��_2`��a^8��OCf�f������w..���m�� ��2��㋁1�q��_���s蔩m��r^1'��p_K��JѸ�Ͳ�(5�%-K�|4��ʷ���w���:4���h��*[�/�,��2888)
m��/�ĸB���l����l��vvO'R,c-DPb	�Ss��p��>@����f��;��ܽ!;{Is��E���	�OfX�?Y�Ԥ�(�(�F�$4���KpH�����)a�qx�W����R4��~��K^��V�t��=����Z���J_*�z�Vnl�~I��@>���Z˚�����Y��]"E�e-ēx*+Êv�����-[h�b���I]6�Q�z��.�����ըOd)�ܓ�����I�^�v��x�X2���Y��]rNO�$fCF'�z��Tv[���������X�5㯦!���7g���j+��ۢEl. '+����S�����w�����A
���g�I��fvS���3y�^&�����!)�p��<u����I�b�,��{�����S/'4s�^�}�`�^����d������N���㷣��w�U2a�/��팴�vTp�D4�~\�c�7i���l������F?�@g����mZBbE�?ʤIm��҇�H{��p�V!p�Z<v�$����u��9 �p�v�4ر�SPȉ�N��Q�q�k�����&;%w���o ��@x��{+/S*���3߅�'&-���b�`�`���S�`µ� �--���K���e^"���b9�{�+GѺ#<C�K��!������-α�+��E��$~'e�����j��	��/����k�se	F*�!��l�R.Sܥ zPj�:6�����&'۶�1�`h>����o�B��.�qu���H0'�V2���s9̃���w�8m�~Fg�6�TD̯c��I$����o18l��r��!Af���9i����G���
�1�[��N�X-Z0`Ȳ�(፛�t;���㧴��'��X� 2%$r-�F����b��^̸\����]���I&ҫѲo�q�)LYh =>���3��2t�S�����|�9��r\�e��x#\r�6g(]Q���P=�%Ӄ�g�5lΘD�֯Z:����}NY`mPP,tS��*?r�L7��9��ԟ��wZ��X�
5 ���ϙ;�2A`G����<թr����j��j��O���P�t8�!U�9��oH��`�V�ci�a�� Chɾ�l��\�}4��fg��S��>�Ƙ�G����-c8OR���{�=��cC�f���V
��K��=~��t��r���0-{Û>IP�E�vx"^I�>suMzq5޴�2��ڜ��m��t��w�o��P7:�7��c�	f�5�C%�v��kY@ǖ3�f�ss��B8�u�ӕ�}������x���a��?S�t�hil���ĉa��w�= ?�O��P)I�X�LFh��pf�j4��Mf8�Q�M>zK^�x����P¿7k�2�:W�sh�|>u�+�JpD��$�1���r����v����9܈FhU�
����ъKW�%^(at�_�H�����%~�����z���b[lˊO�H�L֔&V���X���	���rDȖq�&�}b�ew���O�ЉTf�yd�a��5U�'�T�����V�u?=���q-RX��`͖����3�®��8�5u+Nj.�>�Фp��}f�=Н�lF$T�y�����6-c=��\tc(�	\�K�@@�Ҽl��Y�3:�pU�fK�;)PA>�?��x�d-��ސ:�A^����Qlk<�[��#l2�ڭ�g�5 x�7����啲�X6N�8uD~%$1�'�]RI�����
2���.��L�SIX�Cb6��'h4 ��bp�,�lR�p�_�*Ή#�.����\6|��+�Q��S��,���;)��>����HV�ef��x�Ͼ���S��d�d�#�dRS�Cp�C[�7�����`�RR�d����S���_���Dɞ��:�d[�uNg���@�/�M)��w�Tr�W�'C��|�^�������QTG�y�֝��f�iZ�o������x�w^��{�i��Hy;�����
��h�p����7��g90��r �����q`A@UZ��0�9kb(�2�V�6��pQ��Y:W܌S$2���ie���
���F� ��Ŕ���ڙ�V`;�N��_0�iv)$������8�@~�1�e$�#��&�����l:��Uן�ٚ#���5��l5줈���a�lzp���n1�B��z������7*d�vZ�-[t7 �����~��oM������S���}�9ǃ�tU�M����y�/���羦��Dx����8���<`n#��ѼL���;��A�����!�SX�kK�D��S�X��J1����Kv�k�u��M�=�ҳ�����~���e���Q�T0����u�5�AK"���^��z2{&�X =>ݜ�;�`��w�s��M5H��a�}@�ˌ������M3F+�>l4��d�+y#8g���mW�3��`���@0Y1j^�M�9�|�n��$��JoY����L��P)#�����s@��D�(a��;����9	/��ps�����-$q�|X��H�F�_�+jr&9t���Ƣ`>�w�Yr��=��l�V��ճ$HR���a�=�ݹ�M����j�F[�Ȭ�]� ���<�1��WJbo�<��/�g��Z���=�=��y�r��{t�Nfqw�H�����Ϲ�uo�D���TJ �UG?-�L��Ӻ�[a�d�Q*ƿ�^�t$�9�V���/�0k��>�ļjN>�e�0(oN�{�*�hI��wہ62?��Ѧ�.{��Q��m��Y�Mi'��ij���!���m�f�ZD�@�S^�m
|�Sd�Bi��j�ѥJ�q�9���8�k�F��Q`���DSA����=�PU�d��B����������"�7_s�}N	X@L�f��to��/����Cc�@L��BJ|���^Īq[>��v����\6��!}�l�+�PP�n�>��O���1h��iy��2��1z��U�a�di)����&^B]zX ��#�s�-�A2�	��X���'�r��]0M:����C���	�b�yQ[�%H;��N�A�G�%��8a�u�`��r�e@�H��%лA�������F-ԛר�<b�����ˋ���8t�V_���Ws�PLWPݖ߶�����ym�����f��`�" ��칓�
�τ>�y��X���א�t.,<B5<Md��� �yl���4�� ��-,�+ҕ�2��J�{���gs�b�\�~���Fl�Y�ڭiko,J���:#���6"-l���7^Y)��O�B�W#�.!����� �A�n�b���*Z���A�r&}�Y��n�H�ۻ6�C�5��ڌr�b�-�YͧyG�.@=M%�� �Օ
m��Թ��ϝ�B�N ��Q}%�ie���Q� �3"J��k(ς��U��z�� }8�O����T�`������~�������*���t�y+����A~�[�n�/BMP�̞���u_?���=���M]�.!���7�>���G����rR͙��
¨"�l�=����n	m,����y:XHJK-V5��Ux
RBE 6#~���������'��,�}Ӂ� ��>��v�:s�y��=M�I܇���c#JÛ�U�cP�[��8��z��6iL�i:PV_~W�"�9z��ꭹA��mD��9�/�v_tOdYi�=�������BPCW�������Ts�e����a$po^]����`��!\��J�.f�,�p�c�����F�_�C��5�sM�y=vd/W6x�V8KL"P�/�e�c���_g�H�:M%Wb"��@��@ٓW�)2֟b �F���x$��-6���u����'�l��Is� �:��:�a�Cjs}щ��:��~�I"�����^�l[|:"_m����&7k h�#RF�s8Mn\�(��A����n^�R��
�4�5�2�gV���e���t�#�R�{ç�B���.�#����-X���� q|
�^�h�����c��cg�C�H>�L���,�(� �e	5ݏ�2���a
����B4�u�C��w�B��1�b�C�V���m����Fnd�v�"mzFB�����O�9|Ҝ+�_�{��%�UˆBl��K��%d��Ř�ʹ\>�0���p��:Q#� aԒӧ���	��'�����aLz�]١�!v�b�e�}O��֧K^_by0��;J���~(�!k5Y����F�]��$$��>3��bS����A���������Ђ��Bz	�+q&����C�XJ� 35٠�9A�SGw�*����
���{28���{�w.p�o�^�$�'�]ʇ��B����3B�64�B C�K�<6Pc�B	Bs�Lm����K\͎!�.ؘL�І�*�{{��<�#wgr��#ʚ�K�_n�m<�s�3e��s[�"s&����7��+6�B�c+q������L��:� �>�V?����c_�l����Ě��5�m��z]+�U�?����ô�&壾�Υu\Ft/�	�?}KV������Jr���b�,�������y|)6�o�w^f�`n��6X饴����_�W�'�8�F��������rH�&y��u��(p��%c�Dl���V�{��1��VVbȞ.�~�識T�ܕ���	NE��\�#�:�N"�Y�J7`����q2}�C �<����H�s�?����j�*�	W2�۠��Z�d����2���k��{0ґ�[V<�*���N�Q�< �.H�!�=Δ�KROX��8{f2E.�H��fÖP�A�B�k��/\���p)�@�#��E� �wp�.1��� 4�=��,p�7��5�6�F+�Ԕ�L:��6�j2ͤ>�0%�W[z�������p˹�xD�
�F����|������e5��X�-6#Xh�]�>mי���֓b�e��-Ʒ����ң�C2�`�}ɢ�J�q�eO�%�T#7�ԡ+�E��*��Z��q�'�ތւ����k#]����˻�ӏ/�,�Z���@�-�ER&��1YX46أ����*� �Q��ŵHY4��C�����BsNj���{9b�W0�:�B(i���x�E-�|�^]�,�՘F[�u���T�3�O%��_��1�R��5+pH�Xm��^\��P�R��z2e�_�z����� �I�^ݒ���ާ*ֲ�d"Y�������L��?-_�.[(}y�\ք��/���:<��%a&� }�:���)'c+��S�h���ڹ�ʀ���||���Z6���3�4#���{:�~}��ݣb`Nĸ��6)zz6Gɣ�PS쎡��RY��
,��8p�$�����y ��b�g����/HB����֠���}Z�WE��(<]�ҋ��x����<�Y[���{����%�pP����eZ&Q�rj�n!�#��6�^�>���_@�7�`���1\�����6�m���������&��. �=�i3a�	�VQ:/�o�����qcS�,�I��)x�T��D窮�yN�ͥd����.�3��i�lf��q�X�>u���Z��2w{Ҕ}��4T�*����;��*���U�~�^?�|3k�5�&󑝌O��=^����|�x�I�'U׼��TxG�����"
�U��k�ɥ8d~_OƮ�d�`H�da�I�\Pp��gtk +0����<���Z
]��A-�U������k�d�^�uڲ��v�̭A�g���\�j���E���~u��R>������Hpw�
�Dsj�߉K�Yʟ�y=��ϣbL��]�lGM�8���� �cd���OJ?xi�xs��nU���4��/���������E�$����֐����T^9�b@$K4��,9E�Sr��=����TÎX����j�/%�8R����CG��%��x5��G�z�Y!e��͉�3��O9�@g4⼣�	���faa�8��F�� 6B�(&�*�!�V4W
���a.�$�4|tkL�4�_I;����44��<�c�^��t�1��$'
u�H�q#I����ɧE?@�f:�����O�ࢱ	ïi2��{�&SR�#�e�x�s��J*)�'IB@�8�Q@y�F���(���a��G�0��$��0pq:�<�ٿ��}a1�r���ѧ`=K.�b��nJ�U��z1ugڻ�Q�ꭈ� #p2��B�+�.\:z\W�O�^�S)Z�����a�/)kj��k$zw�� ��_��y��:S!U�"E��Z�L�ЄMê���)y�H*Kƽ��u�;ޑ���H�F��B�d(���D��:��)8Σ�� f["�?�7z+<c��ܟ��qR��?@��rV��G�)������Nf� �{��4N-����\�-�D�X�ѳ�5�@�j�h�@��{�vu^��i���S����OS�h�
*$E�Z:
Bim�|'�'UBwh�I8��c�F�P�e��<ʲ�o��]�+C���� t�S'>2�S��Y�4?G:"�k|S�^���*THc�["�k:P���8���0�$�Ѥ����ag��!~��m��2R@\�B��+�N'���.@�7 ������v�T�%�*�~.̎{���h��r�;֘�Cn�,bnǋ�4���$@0�'�R�D��U���@�>��'>��Q�7x�~�o�6�Wc�����)��@�,>�XG0/]�ض��$�z���Z�Qe�+�ZP	3ڠ�a�އ�z3��m=�ľ��9k�K֭{h]ZM���k!��W�E��]�AS� �J2�u���ި"�w�c"�����;ЬKB�N9�� DN�6�z�|U�5u���>�[2��Z��gj�?"�`�_(����@��͏������P`w:�����v��܂�/�S0J�O��D}�=��l��V�Ӫ�ՠf=i��X��(��&��.�/���QG�"t�X�U��ˣ�m3� \�z"�N�j�Ѵa�4Ά{������wY�GG�(oV���d��	���6�J.#�V�su��"=�- WUe�����vcyl� ��Z>�5��y��X��m2�;���+�׵ׁ�������Geu���[�����L�onu�h!�+�[B;I�����3
��F�A k����J�s�q�ڵ����^������Ga�����yx�8��s|�g"s��!+�����5��I.���@@��4W����X]߷=�{BQ�|�����z���kzB�Zw�+�.x��m��v���%/v��'��o�?�r�u��c�Q�!�TT 7擺��rb��� kY������/�7QuG=�x�1�p	�D?ހ��}w���iR<��/���վ?��nP��J�Q⹡�=��O�Bᨾ�=
k�����,e�?�0��
M_J��y퀹b�Iy��GH	��I�4��:PT9t?���S�T�!k���U>��̪����%��X���� x*�SG��X�PIwt𶽰Hw�V���nQW�0W�������d �}���<FqT,�@�]w��\�R��IAʻd�[8Z�g@sCI���3��T��+��Q(�j|ۍ���K��(z(�!�
��y��då���� Q�_�Y%��}��P���������a��u��[1C�:?J��f`�Y�˷�W/+>#+��4����	��a����tz#ܶUM��WOhW�۳Hጿ�N�6�\cAݏ�ڈ�JCf��f�G��v�򎥸��|;冁��{ڞz�Cv�'��\�x4T���D~�I�\�@���Ӓnó)��H��*D�"͑��V���d��5' �qP7cYQ��Wg��pP�`&#����_%"�J��.��r���{Ӫհ�Ȅ<���G�����
��ۥ^N,I�m�{���8��m�vlg�؎��o"m���U(�֯(v���/u�+���q.� Dԥ� ���ʃ�ي�:]�vtn�ҹ�΅˅��@�'wP�� �w�b��rW�?�C@Uԛ���S!��ZA��Mޑ1�\S�r�	�:߃��J]��՚�@gB��F�5���xb����<�ar��xh�ۣ3~��G�: ��CG1h^�A�G���xn�?�kG�a�����s>k H�(�h�8iV6[�}��dh�l�@�8M��aQ�^�(ޢ��ц�子Q�9������i�mm�%��F╂t�8��A7Ħ6|'-�#���=��Π/K&�^wt��d��5�#�ԱrI�R��Ǿ���W��!� �����O���eDdkws��w:N�{��������)�AM�t�nl]ڿ���.����مa�h%���>7��Vd��K�ɚ.���J������u�O��������L�P����sҵ��Q��V"0r�?�f����?#�~�",�G���y;h'cR��a��m�^{��7_�z�e���I�y�����P#���\�Z�C���)�,O��P�����Ò�+K����h�Ǧ`*�C�-w��8k��{�øST�i��,^5>$�d=Y��'�
3�g~� 9_i�P8�+�P����'�Q�#����3�t�D'��ԥ�uu^8��CK|2Y�j�{\�����S]�_x�m���-kl��a����`�GAam%�)ͦj���9/�%u�1 ��W�+��<��F�u��s+�[d��⧣qK�zj��Y� �:.�ݍ�1��9����+i0g^H��~��/q]�ǣp/�?�e���fR$�H%�L��b5����Đ�1d<&T �`
	��ȅ��f;�u�(Y�b�G �=i]���G�'\��V�v?6F�����LC3�eޫs/�*x����u/u��q����R�0Gl���m
����[�o���J������OF��?㉞
t-[>�i�<Qo&&����qL�x�Up��lC�8А�`�_EVQ��f�bR��R�r���ev��z�v�̩��1�#}�lPi�5�<,����PEQ)�A�ֹ�z�Ic4��)E[�9pҺ�l��;�D�����Ꞻ\L�\��n�
d��S����Px��"1���Ө��L��j�A�Gt���M�r�
���V����n=�ު�#���g�x�&�?{��ƟȢA�l�'u�o7�{?,�>2��0WX���H�}�[�3�Z�����
�w�x1�s<�<-%�	qk������ZvX���" K�0A�E	����s��aA���� �]�8;l�ZE�mf�
ɭG3e*˿���SP�#`Ƅ�E&;8����uzت<�5�Ӡ��/�eƞ���%>��(o��N�!I��F%9�����K�kV�Z<�.��_�ς��М�e-��c��]Di�������G���y�Q *��&�j2��gM:������Bq���CH^�X��|V[D�(i��ad�ky����+t����%���\)��<��;v�Y
��(ٞl`�Dj��"* Y;X���I����s<[�aN�o/�	@(�����H�������z=	GRT���v��G�dh�]�Iy��nV���2H_�O��e.z��UegpisL����[?s�rH	Ϻ�t������>������YY�y,�$ ��J@��������>"�y����h�qێ��b>D��W#z�0��'���vr�RΣћ���ET:�%/�6�E��?�c��0�[���>F;��ߥՎ�wl�j���Y��n�����N��p;\]�љ(��m��j���΀�\��{@)Eb[�-5�|���R�d�ʌ_�"�f�N�LhE�Ґ�u��(Zʿ.�J\�W79��w�#D����m �$���,5��U�*�)�9���Jux��}�W=���=:�6�`� �0�%0+�d��I����f�o��{�^Ħ����f\kpd2`�-*��U�Y�&���EQlQ�O�����R
w�"��ƃ�5q��	�4�WAy��N�vj��_�w�~y��`�k��=pD��a���G�� �ExCI�dc����ˢ��A���� ��X���' ��]���q�����������}��9�<h�M.�� W�P�VyK�98�A���	��_>�$��k�6��~��	~�K"IG�U����X�^.���,�P)*sz��S�J%��Ap�^��}�����W1�$Ͼr&&,$~�SQs_Ң�k�ɚs0�u�!�)���c�x2�$���\J�Ci��������v���r�;T�aН��b\=����7un���	���,��:H �<o�M?�h)�#�Ә�c�ձ�-ymZ���
Ձ��Ј��_ep'���f_�S�d���BaE)-u�B�YN�V���o��-�s\��i�����v�I��zVd%�~�-s�r���u�a��۞jT���2�.������̨5I~�/��8:���y0N��\Sq�^�"��mT'�����gG���hR���wP!"#�Ñ����V�0m
�ɶ︊@�j,��;蠮ÁD���щ�]{��	��%�@�c/���%�Ӽ'hoq�N�UC)�(:��rBH���8�ɟ�/>k� �b�7��c�%J�z(" �vsAW�z�p�\5zj��iJ��c��2�D^&1�SJ@&\����aI�Lb��r��x;���.��Z�_>��cwz%HIv�s8�yʅ�{��b�݋�aNl9#$�@!��|�)���R�8��;��"�7ņ�D��[�k��/V>�"]�M�*$�ҳ��4�r���U��{۴����Ј��Sc������|\��R�!�:�e��ױ&
�Hh[��\�����OR�8l?�yJ<S�8��~��8�'H��Ǖ<P{9�|l6��4�P/P]��x��.v��Wz4|΀�n�[�
i}�����.A��C�h8���.��^[3�L9V����?N-hf��[ I=1�W _�� ������f
����B�~�����H	L�E/�3H�Z�i�C����%�K�%�м�:�P��b��k�<��V�&����}�.�j��BCѵ6������4�6d)h��R�[�I*���PB{`8�ʘ�H���o��P�=�Ϸ��Ϸ��q��#��f�}��q��r�86�j��wTQ'��у=���am5dڲ�5Q{|�֙=a�:1bll�Z�|�7Jy/g�
�0v�R�K��	'2�b��z$��D���
���c���QW0Rc����W�o�4�>WDH���;���1Z����< �f �������RLyW
y4�����uT�>�[���;S��:qb#4�C��X��"�>ݒ_�i)��PU�N�(x0,6��X�>���[�"��%���H�a]%'�M����;\��<��kB�����L	x�wKt��S�e@n�ʹ��xf�R�jda[�C�D�"�ϭ6�r��L �`!2w�O��=(���|���L��ƞ��[f�.���F�>e�ׄ<���?�L|��Ϙ[hK�pz�ђ_�4��<E��T�Z�ɛ�%��RA��D�����%���+I�r{LL�9���
���/�?T�l~u6�+hPh��5(�qh&YcG�{7������oe;c���f	d|y���r��q��#�<�����_�\ӗƺ�H��WC�
� ��"Kp��l�cI�穒����:W7u�)����hmf��
��k#��`��Q�M��n��b���+�HXt�Ciw�$�j��]�W����&� �d�e�7EG���t�?�P����o#���<��s{L��'.��[#=Ԫ������@����0�#�\�X:�P��	��*� �.:��	�9��(�/ɗ�1|��$`M�_���2�k�?N�����:c��_k{�~��T�͙j�>�]z⸞N�s3'�"r���b5n٨v�_�hl��k�Y��ƀ�2�WR�� W$�mF+;�\Ŏn�^ݤ�HtVKm�v�H�
TP���6���P���F���f��;e���ŮB�[�G���zm�i^�U�A��&��ώl�G��8��ûxKw>+ԯt�d\�:98�"x(�m5Q��d9���c��ї�0����?ه��4CL1��QXq�Ҷ�Ĳ�%m��ß���Ŀ]����Rp�DW)ˣ�_��O�N�aE>'M�l�x�fbs�Cp;,{�����T��_$J�Ojt��wZ�b��|����9��G�%�ї��eM3����8�'cvЌH�X�J:�lV[z�fE���FO=I,뷮MԚ��p��)V����&A]z�L�_�.��sF�D��`,n� ���,��*/��Ez��Z�j�vߜJ�{ۡ�3�.���XRe�IP������[3�tuܚ^��Y(�h5��w���҇�H�(�<��w�"j�sY���$߷��cd��:�(�˟E�|Q������� '�-B��;�	�����.����{��7���_��;��n�=Ԧ6$�աh�mF����rF��?�����Y�%�?Ѱ����D�����h(���+��z�
��vJþi�ìQ�v�@�ƴ�6)�2#��]��%^����j}�TwQj���2ڠ;���r�wbཷ���_�s�ߧe#��;�x2é¥6ժs�h��3��liQ�d�������;���/�����kC3���Xw�WU���Y�.����u6Sq�J�k�YF�k.Gq���� k��黪�����8�
2���7�/h�KN�s�4L#$�e8:��$��{x��.h��ˁQ�� 3^�?��>�-Dp��|�=t�\h/�3��q,������"�s�hK��]�*�z�WAG�=d���Ξ@}��fh>ͩ:���;َ��[�x˾��m��v���,��m <P1��c��5�y�Rjp5O�=��{�gwz��˅�D�{����H������ܐ  ^�-���&�?���k�8���P� s&��v�+1��R%�����kaF�}?�)�lH��(��Q��wc�dҶ�*�{���O�c�U'1�i&��[�k������V޵MR(��n�ד������5�c����7��q��{n��lq���
{=Hy�|�d2F
V���5+��7精-S�y�y�A�1C@��`F�g ��(�Z�\:��g�<gDc~[��f�u�H2�(	'�Z�o��S%�V��g���f�75nE�	:u��Pf3�U!bjU
����wV�!k�H��`�AZ�O�o<+��ćK8����Eݓ[*NCi�N���:��*�-Bk*rb�]����9z�%�a�u�g�"�ˋ���GGWA�>��:y���{Is�C�RT�O�Qr��]��46��;��b�ď��&E�<���s���oW�&��r��'?|;�7�˦��S��ʜ
F)j�~Um�y��8g���J(�Ҿ#��&;�u.�MԀ�3Y4a� �qlT0B��������`� �z~�ɇR�����A*A�t�8D�gFx�`Y�}�B�Q @�� A��x�uinN�Q���gź�|NiQ5�n�fIC&��C�߭ �ԩ�r��B����S'|�����>qN���$�]%�Z��A~k��kO�lԇ��
E�[Q��9F	�L�)SM���<�2"�@�s#rD+���?X�%3t����2��@1/R���T�,�G����6�w�9m�K�r��]'����2�>�]�}�#M�R㸖hH47����	�����~�O3�q>�rytw�&�Hژ'��r�>�8�s�_�嵲�	X=��K�r��r�@�	�ѿ���*2�&h�_$�r`�>�F��m�t�~Pm��!��o"����F���?����\�q���ʁ�hs�F˩C`AB6��I�<9]z��W15>z����	��g���-��3@}_xp�n�}��.��l�.	����"7�B�qk� [s����x͈�o*�Џ��ѭ���DgN'-;�(h	��}c��𣯳b�E��A^V�3����]�3���1�X��O��YٗJ*S�Y����n�W������V�xHe� �9z�&'�r�L��g=�#�Q�o��$x���$�՛�]j�h�>saf�Y ��D�6P��|_�o��-�� OheTW��.#�K��D�l�u�~K�gE��C{�/��'�$0�ԺJ��p�v/�ԀWm���a�'���ӗ�sZ�lSv��|8�ݘMz	 ���2��S��iqH��/��O;L��[�ł�1Q�/Fe��[�uru�
�L������q���X�[�A#���SҀh����NOV5H�x��j��_��Ž{�>�{Cr�h4��H&8]���In�H���������tn;�	���D%�r���O�[��(��?�?�W_��-I�G0@��F�d�U����R�/�r��*�f��<���Mtg�+�CB�=�Y!��T��0�k�t,)����oqt��u����%��&���	����|�QiC�YCO����ڙ��sM�g�vx�J	�S�;/΄����[X����(�.�#�����Q��[,�ԇ��_�˕3ᄲ�p�S��������a�H��#3��|�KJ�W�._�U����/\�� P�|h�w/ݥWV��2�uT��D�`8*$7���s�a��;:�f��nQF��/�� Xk�([a�O�kg�}0�G��gP�������g��߬����v���J�Q��ΰ�;)q��T_m�'��oZ=�ߥm�1H+��X'��Ԫ�������Jt0^�ʂt�m���RV"��[��� �����$8υ�������%9��A���䶖OI%��;�j��ׅjJ�l��C}p۵�K���R���D��e������������ �t��Y2A�﫻��ȳ�����ж�R���Ě�:`	*���CV!���]����.�1�����n������L�\`J��H�i�	��f����8E�3�S ���h��3�.mj��][S��k6�:��đ�/&��S�Qͥ�Z����a�'O�XM�bC
0W�QQ���=�+A��U�S�r��ݞ�{����r�����Ѡq˩$!8��=�����3dJ����P$�Jg���J�%�abG�|��A�=!ИfH�.<�겖�Ɣ]�]{ݎٜ��� ���v9֫S%�0-�9�	0?�c�6��^�\\�2�Y�󜷑��B��:��/�@l#Q�iV�D�:W}K�g�]�+~�#N-�Ubދ�>v[K��� ���Wr��l%0}��%!b��A�Z"i��|��W�x��*�T��h�t��cxo�d�h38�ܟW�g�$QvT�"�;�Ӎ6�B�0
��)J%.���	�4�]eV��kp>qZxZ�9*�_��CSHB�ҋ֌�L�ĩP����B�q�l�?��HC����^��KR�[a�h:8>����Q��fsz�(�aɸ�6�$�,��g���\#�c�����z��T�6@�\�ݠ���'��><1�+r�Znҙ���������x(
.x�Qo&�U���ƻ*�7�H�J6��L	Y�����?W�mҶ�%���F>9(!���X�!olqX[B���qoK�]���TY]C��\�SJ4��{�S
<�"�����^_T��L�Gu��}M��iR�h�2sh?����f�vvbz柂�pz��h���-���J��eV.A+1�[8���h�\��r����٠��ydHK>r��b�g���c��E1�����á�����i*P�c�q);�<���n��vn�/#UUR{'�,�cz�O��
�'x�D���f�y gF�XL���E� ��=ߵ-l��C�D8�^���?����NM������Q�H �{�c�N�B<C3���5�>��zYi��!�垰��<<�����V�2Cc�"NRՏ�y�1)��^��a��³ޜ"c��
�%���N� u��0\\�W��[d��y�BP=R�PGً9���)?S��Lb@r�W�'UcǇW��0� ]�#��n�~�< ����Qt��+eBje�q5��s¦K��aB�'�*6 ߍ�X9�*��z%�y�c`;��;��L����&�Mħ����H�'����Q6(Iv$ϰ�M�QC�sVL����tw�Q0I�	��`�;k�v�"��C�)#9���yV]ݩ��>��\~�8��k�g�<�iؖ}�Yu�3��0A��YPh�s���ڤ�t�oW��X�A,N�tXD��O���&�Տ�Nѡ�G	'�@7�����i/[%7���L5 LI�L R$P��!m��V��9�5A��s�fwb0&�� W��[�,�k����Z�I��g�Y����6����L��$�m���aS��UN݌����o;��fsTOu��=n �	��Tn�������N���p������/�V�V�|5�O.�.�{�@R�5�iĖ�At>�k���"��}e��+/�f�	pt�!��[�:���+m�8粆˸n)S��n:C������HqҰ�!0�����b��Vy���h��n0�Z�k���I$w�"�u��?~�������b��]�Qa��k�{C*�:��Z�0���FB�O���G�����x��d�)	�K��qpf�b:˥\�k�K��eT?��@��$�[���3>lD�
e(�k��ڳ{�*tn��oy�O{�_	����!�&�l�-�:|�ҿ�_��d�`�|c WFt�fw63n$iq�]�қ��lљ�IB$��d������G�B�J;ߴ�}yDS�}Ɨ�8�.��]����_	�$�Av��Ly�9�qHE7�}O	�>&}{����@�9���,m@����+h���]T�gT8�Vi��`��ٚ�ّJ$��DҫJ����:�4h�Y���c%�˵��ŵ����H�~;l�S�7�b�5�'J�TlޫC�Y��!�Z⼪n��l��+�4 �a>UlE�y[N
)� d����[���qQ�����������烝��y�T)�̞���m ��`�A�1�ԧᜉ̭��E3_���Fw Qm����A�b(TL
k���� ۸�z������#�u	�6 ��U+�</��������`,�1L���N���0��u�w�7��[�p��>پS!LLA�����Q+�M��ߓ���Чg#��{�Oڅ���{�i��c\_�0G@	�D C�&��bPS��@]�x����Q�'�eml�g�@r¤^fR����F���kzǒl%�kC��Cm�����?L���i�Z1�ů�*��1F� �$}���"}�_�����r�Wi=eXPPX;��D���ck+&�i�ZL1{��h*����3� �47���Dˆ�{�YF�Oe' �~���%eU��-�9�߄�n���X�S�r���߃뻽�����݁���V�h�#��!�ݹ(q2ä,�}��_ �nWg���"�sd�=�����{���3���<p���D_��8�*`�-��wt�?���y�J! ���;�,U	��Sw��{$��tq�6�Pm�h�yBo1c�O׵9����hаM)�t�N�T���(Mdm�\0��p�9��O�So2��9I%���$�]�0JE�(!mɉы~3ƿ�� 7^/ �В����s��R;�&�+	�L*h�Lͤ�
+JU�����"��s�H�s������\�\��|�tk>�J_k����TZ�<Ʋ�9[�@�跀J�1��;~H��[6y
ڶ^����O56�ýշ�M����X�O�6���&�q8�\�p[y��hs\u�{��q"*|r��P��tgd���!���3��)���C��� �����<,�aR��^���}���6؊�aN��z\uA��0�MPb�R/�E�X�B���,{]姬�/ƮEX��!���%2�h�+[нt>�D�����A���\��w�V#*bST�y�?�Ӻ)<�H�J����|8��LQ] �a��qQG�̪<t�����*0�)!uT��|9�h�K���j#H�<9<�1zKD>���^�wj�n��a��L�t!%M�?������#i�nug�Y/���T�2c]��{o�^W�Eg�,�-��.}������(w��!��Ȁ����JVA�қ��������<�_�P�40l�3�Q���vWut�3��x�ND���2�D����j��0Y��e��@-���GY���"�3E��1��#��*XN�3���%��!��<ĥ9ۊD�ߘ$�Ivs�Ԑ���~���Z�9^�w�ŽW��
L���G�8��s>��xٴ��7���du������ ȯ�#轢c��%�]x"�y�D
(��8W>RV�5 D��X��#��WE���y��z��AP�]X]�&i`��6H��U�U?��I@�lp��
���� �|_�"�-������Z}9Ɋ*�f�H���^����$��[4<���`D�ݣ9�*	$�o��q����Bz�Lka�L�\��h��#�=�Q�cI��Q�2[flE��2��7�Ғ8<�G��,OFwҲ���qQ"�����@��
!�A�[��5;g���+t��#A�/�#���-������iah�����ςl?�+[�m@�lCs@�T�A�)�-�*�!c�Y��}
�m�2A0vP�
"�<Z�t���ǣ�@�ryq=�2H��o�j�`��z��|�7Bxݱ��(4���g~�\����h��F���/ |�6̏�����+ǥ�.U��ư� D+]<�۳;�(٥�z�����+Ƀ����@>�ǀ���ոF�Z�����t�M���dCڗnw�Pm������4NR/�^";��2r�L\R�C{�R���
�:�F���#�b��d��t�8�+/��-����o\G��+��%A ���^6�G�*H��lI�:ܟ�&�� ��vr�����8���ȱt�"q�l0��=�5�<Ͷ_�l����ہ�sID�i����/>V��c��E���_������Vp��{~K2}�ĕ�y^zS���-�S2*dOC���o�Vp���b#�}���'�	�+c*}WѺI��<�/GF{̎��gܬE0sU�l��1�1l��u�PF��Q͇�؆�f�D>
Z $8-_*�lf�9�1�pyo�ө��L��=O�?p�[.�2yv�W��N�f�J���/q�9J6���O����+z�{�P[*���x����H�7#.��۪C��-ث4Ti�Ԏ��A��e��X��n�IXI�)�K�#9����|�8<���������s2^>�&�[�#v�J<��K,~2������wB�A���<��3���z��(|���Od��̷�۴�=��Y0ګy�_�� �l�`�n0�vd%��蓉^w�L��"3=׾��_@Cf��k���Ϟe�Mv)�%���h�{My�]���u��<�(ģg�y'(ޚp�Ҡ��0�wN6]٬ϗ�z��(T�d���@�A�tW��n������2S;�c�E	`Y  ~:���lH���z��.3v�X��"� �d�xL�n�|�܀��^�P���ꗰ�N;�>o9.���댦;��D�3�i
H]zR��Q܋a�xU�[��`0*�9G�&���
��m޾3l�\��jV�I�A㳁d��Q�?�/
���Vkf"j6�erW$�qs�ւS�٠#�ywQ�͜ �"hp�qܐ������R���u�v�2�&7UJ�K1�f]uv�
�b[��Q���r� �I%�h6x��	��  �@v�S{SQg���qvWOB��婠�-X�0��&wy��O�]xh��j���Z�ZK��eZ���>�yl&9����Q���|�.e�b����k��Y?�|� ���sTSǵ�\��@m��碔<�|���9a�MF�0ݨV*h8�e �AfF��cvh����b�
F�zjAQ�UG��Ԁ�+r�k�3�՛ᅡ�y��b�����$TM�tCDaٱ/��7<h�A l�LL
��O��Wi�߷*I�n����E"����<�]}��Xt��J�m��Â�tа�A�CI���U�v��/@畕����ބ��'#\WyH�C����}�~�o�S��&��2J��H�`*V����,c�����|��6<��@[�:D�8��G�� u��b�Cd�5j§��z"ē�Zs.�!��XF���m��l���~�lw�y�AZ�xdo�� /bEnaa�N��d����w�1#
�c�n��Y�w�0O�"��lnXA�߷aw��S��in�+Pn��,� �^\9ȩ�2���iwC���ps!�$u�v)�Wx;=^�����!��I�b���{y\�GG���Z�B�EO �6�ޅK�q��}�Pf��e��J��g&�sZع��m�I�J��0���5�1q���1�QAg �-ļ@�^.6�8��e4�*O<F��qa>�|<3�t�m
�uc �/u�p�к!lp�=� ��
�+�� (�}��d�B�+!W}�*y7�ݎ�ww3B��D��c�+Mwr+�\>��;Ҩ�N@��}��7������T�F?GeY�ŪʥhKp��f��8dBipr�ʪ���񞤺ǳ���M'�3�ړ�t��>k��J��YS߼z�׍��n ��(�ۂ��8C�*��m��vMMYI�u�J����0C�i6!�I���T��eW�R���z��􅮧�9v�����Y�d��eb��99��K�.�cv(�iκ�VU�#6��_f����f�Y��T�DkBwp� |��g{+y:*�P_��Ρ�q�R�0A�������Sa�|�W)�!q	�Pp��-�ܝ���w&�y�u�p+������	�ƃ�j�秩]*��z�T���L�*?ᗩ��q����tVԯ;��)��T����wM��c��k�g V���f���{�UD����l#����Fu��jf eQ~$}�Q	(t�3������p��*v]�Rf(��2I�=l��^�&�1�ӪQ&I�#�:�c��k�c�)�qR�%n�F=�R�
��Q�Ї��_�7��L��s����ھ�X�����e;�}u>���F�:�c��]���>���3\[��	�����gm�)��m^���8cWYd@_���J�U:�S��"�s8�����+�p�J?�gq��%����,�n2x+���N�[�Hes
J�i&>~1���]��\����߯�&�*���fU�S�z��H%݉�,)�>�Y�#ԩ������6{h,�x��51Bv��ȿ<��/��{��v6+�$��|L��\�-�.$RU ��}X��V�&��1S *�/J�'�%d��0�%p)q.�2jN�5��c�u�e�-��J�)�k)4���@�d�@�̋�˾��%�K6���Txl���vPz���p��baBX�=^T�1�(�}HBfH�QV�=LR�����e��1w��a3D�ݥޘY�զ^8��^$a�q�?B�.�g3[�`�;�����6�	ֈ%d��h�+�6�}���1�񡶍��1C1
g����z夙��tm4��M��0�����By��,l	�R�?}���hmad~+�\&�vB�.�����[�C����2{��H�����0�X:���(�G靡++f	�
1`
�-�!כ�8��NcJ){s�i�ʀ���+`4��!i�ؚ,=��6V���^��.��k�l���B���߉�y�O�R:�jy��I^^���� �W�$���Ü����Tb���u�I�x�-Ix&]�P�7���٪��t�x�?����q�(�����>N_�3�d,){ҽ�:z�wČ>���_{���ݼ^�Y����ގ�\�`���FD<�e�L���=g�H$��{�ʹu]����l��F�	�m� �k8]�����_g�f�-�0�6���@���^��w+M}��y���]^Fc��hW��<��-�E���l�Z>�/�<��ѻ����u�����b麟|K0L����:"�
�<�� �������W"��ͩ�0�,V��ʹI����ۊ�c�������Xjv�]�����
����Mõ��S��c��&o�Y�su��EЎ��4.��ݳ[=�5�I�=�� �TM�Dz�>}'�����ӿ�i$pjGB�l���\Ş��tS�������_��m�^O������a連}qWФ)�]3O��v�+OIf��s;�q�!hx��+X
�,�-x%�C��`5=�ԑ4>�Rs�(��ݽe�t����h�,'쎧Gc�[�T���>#X���7��)���g�4MI�Z�u!b�n�c���B�~����.���V���A���Jwx�Ɏ��J���䴶�xMb��Ƒ��g�$���/"��� 4�@��8��R��'�'�K��@p����,�����2�?Q~�]��p�5L��ÑD��|����;�O�����U�����T{[�D5�b!�d�}���u9uC�Pe$�y2S[�95���R�i�#OjT�!�MyJ)FY}Ârb֮b=򸸥P�E@��c�Ge�
l�qߵ���II��7S�K�#�.U�_rɢf�q�4�w�q�㯣��a1	��L+�h�o��8%��jiϰ����j���U��W�ˏ4E�#�Kxt��u_v��o�3B^Q����O�s>�7���!��&���3ٓ/׾��M^���.X	r��U��ۈ^�5�!I�ubm[����?��`@��?,L``�D>��\`��FR$3Kӷ(�aqz����J ���:��$V"5Q��!vK(�����u���y�z�ٌ��Y�H�S�A��X  �몐�ʧ{G�_!:��� �(�\�Ky4��yk��cK��j�m@���#�~�~H���J>`m2�u��.#K�}��voYzɇ�+!O��tH[��M��Qg*}������]���z��z�D�����NM�"dй�/�{<~��2H��y�������|�9hJ��I���Q�쵘��b��.�M�<��H=��P�$����wD�5@$��L���4�Q<��Q?b��~���|�2�Ҭp��}��A�v8���(��s�D���*\��#3��A�����&����s��I�w`B��֘�&+�`>X�IA���Y����[R��_�Y���A�݈��Ml��$��h ��[}������@��㱉��&n� ���io�\"��h�p�מr�g��\-3�v��o�G
��1!Ԋm�)���9��+m��U<B����H����6zB|��x�1+�����������D��Ed��G�Pz%#��t6��/t]��PK�H���:��F��>V���З��\E����+�8�ђ�Z�C��/���������)���l�ؐ���j)���l��¼+��7���_5%6f�{��_���WI�����>�ޒ_��XMO��ykB�J()�	��{VXʯX.`+�����=���p i���Nq=D"d~`NP��L+G�6EEϞ2N��O
PZ| HW���r�xy�f��d��̩Ồxu$ҁَ)!�Q�c�n�l�wK��*Qw���������O�Q!�s�B#ݶM��Y���<I2���o;���������ĥ���fK�U�í�K~�}
]��.?��*�o��*��o����yLAm�F����|��S��ڬ���!��U��<�;�,�n
@�tw�?�⁀�I�N�����v�l�`���D��-e�rrt�S �=�i�D��,@SE��(��[�W�ف�����N-�v=9s��9���;���`�;?<�X4��G*g�D�b�'�O�cmz^�2V�e�S��R<���>��ry��/'����h����T=fN�J����ZH���i�
�`|bP�f�d�t��g,w�m�����	U|���k&��3H�9����d�h�&�k�m�Ϯ����fm|����Z�ס5=f�t�k�8W�Iw�$U!UE1+���tQ��M��G������As�4�S%_C䀾���E����Y@�\�o���{�*uF:a��&:���n)R�2��Dē{���LY0�O����B��y1�FOL�O�ɮ��N;��O�,�E����e-��G
0�o��Jl�"�w_K���k�7�h(XƖW| :<6��iߕV=e���>ߛ1� (���D��=V" ּO�2� �u�X��}$WVI)`:Ҁ�X|}U`�:�˒P"B���i��l����C&wMT"���]�pZ@9��bB����J���9z0o1���ń�i�r��jR�C����ÙWo��i��>/s���������ײHZI!z�Q����ML�>!���u�wJ,�z3@B��d����A1 -�n	�����ᬳ�_����@$5��#�	��rA:��+�.{C?<x6y��"������qP�/Y%K���B�z�@�e��
�KN�?}�V}�3xuٹ�MgX����x�Jf�z�\`3�J�i���۞-U�"����>���� n���|��k�\Ex�[_sJ��t;rլ_й��]���1l'��
Ǐ���1@�)S|�2:�Fި`H�|�'� ���ʈ|���
�65�����&~aQ��8��q��.��*ZT�	-�S�Fy~�1o,B%�Q�@je>��.j��茚�zi�=:�.�_t��%;�������E�L�e��h{5��o��`MG��B�\k��deV�g�P����kN��+(5��S��=9)���fȫc�ӵ>̶-C}h�^�e�6��F�������v���^�q=!�`f�����{,A�w���]4�ʼ�k����0`�T��뮮�� ���}<PeJ` ,�2T!��R���y�������ъ�H�U�S�$���GMn��8^%�^��HJ�O��a�U���A����MB�YPDa��c�وZHKuzX���2�S1=�m������TIK�Y�B����P��U)���*��\��s�!	��sx���?ێ�G'\����TF
5�������0�@=���$	�D�y�P�P�?n�����X��zi{_�`P�%��W�v���4y���uk_�� %�)V���[��6�x���������Y��kE����n��\Pk&(��ҿ{k��X����d�j=nަ�cO�Ԕ��іN���&��m��R�-v�_u�`w��6[3kJ�{�#�;~O��kO�%�=,G���u��B��4;�C�43v��͍�!���L���3��|̣M064V-i\��^�q�,�	��鱏><�M��6�Y@*U`��(�'SZ㇈�e0��v6���MR����ꛟ\&�E~�f=���$��RpL�W68m��g�����-�ٶM
l|ʚ���9�C#��7�W�o����#�ձ�_��kkLβ�6#�r�����S����r���6�oL� �:
�Z"n�:����^e���,��

W�Az���CAR�>�Qnf��y���kz�D���5�4� "'�I�J���=�g}���������z[��DI��P*�N�1G>�'}]�������Rl��H������R �g	��m�sŸ����U0rˢ��d�X&�z��]A�4�T~T$��x$O
�+�\X�! �n����7h�e���2Q��"��t�}ඪ�L���s�R�����^�I���)�8l�l��혙�T7a��S�,C��������&j�y�a�dK����bW;�$��F�[��f�bE�#FD-��6�F��A!K�X�"N��eͣF4��~S�Xs�Z��^��bfabq�3p�����Ž���Է�}���g�`*[�J-�\��9��b^c壝�RRˬ�L��E�18�v��DHU�t���2�uz��r.&������Y�� >{�#�g��\uv�7pHy *��VB��1�����%GZ�ɁRjH^���;�c�U�Y3"�UEu[K�G�7��ze0��;�I	!o$�<]� 	dnȵ�2�Dη���&͖���񆥂�
{O-?Ե_�е����ʤ�H�.�
����rvV�\�Hm�5ύw�盩4�Vs��3�$R���O�g���\ٴ&�KT�z��k	���@��@�+4�JW�_*�/86�DŢ7|D�ȓׇ�J�q��6��F�uliWU��-�(|z@RX���%w�J~�A��� �b��~c�������b�k��u	�?�N��+2�#�&f :@�7֠t���q^���s��,X��_�������.a�^}���+�s���޵J��ԍ�&���ITc0�K0tAz��@�R�F�O����ٸ�1��a饜e
��(d����H.�3t5���g����b�h�[5,��H2a�TJW.�FrT��>�ha�X]�J�]��vRkD�~J`�W5F Z��cq�觻 �n 'O�� �~@wM�؈�*�|]��
��E�X����R ��1� ����Smj�^�R������>^
Z��yX��`V^1[���9`w;��H�9�Zk%�V�tء�%�%`�i��u|F�*8�\�S�Q�c*X֓	��� �r��K�»@�.I�qjxC@��=���Z�F�6�@πIX-�%Q�e�RwȽ�Ll9�����j`�]����6,B[�*�[�^p�� �@��6�������h7��"+�|0	[7;�z�kh�_|fD)���ŧ��l�SR�NC/��[�E<�g{�Z�Ky/Ε>����q���H'?���E�M�p�¬9��_l��h�36G��}��ڠ��
��=b�ơ�W�sm<�p��i�p�hgN�:z;9�e�e�Yܪ�-ɥ<a��?��j�>j���h/+vrX��&�l�d�'a@:%D/|h��ʇk����4!t��3��@�����jˮ�������`��cj�x�wn=V���_;�Di�vϕ���Jm��	�晽zB�*gReFngNJsY�q��d�7��e�K�� �u���*�$jN@~��dHq�!�~dz�ī�@��}8;A"�K,S�I,Ct.ҙj9<�l�y��dU���G�vł�.M9������5�t��5F3�fM�G�봤}�ヸw	���lj�	�곖�mV�������N�o{���)�8'����2x�
�~F1���p߹�Zr,4��q�V��K5z`W����Ǖ��������v�CI��z���Od�ԧ�т3�����{����*��V)וּ�h���J�;��$�dG@�}�-'j����C���j�g�gqaL�+��Jwì4�삇���B縸T��������
@�oW�[����:�8��#dsP�f�şY��p��>�G������}�DΗ��"O�[��i,���{�Э�H�(�:*�F�N�uŮ8���_=�>��j���`����ұ&�#��暟���]��N��Y��D��8
{`�Wq<A,�}�|
��Y9�$���l?D�U�P;NB=��6��%��Q�V���^y�9�A��i�)��_Q� k +v� �kD�����y�e�س�f�'��%>�u���� �J�l񋷰�D�%=�]�ЛG����	���`��,:��S�ä~/6~e���	m��@�2v�FM�̭������@�J����(P�l�J��#WCk)����KCR�)�c�F�k�PpA��;GPt=� �MCF�����!��2������+���ʀ���y�9��ҵ��^/�����<��N̒k�uE��fL>�۝��g�SJ�Jn�DW�A1����8��I��1��,ۂ�1�=瀄�E�^Z��=�`\�Z�ɑ�<���>U+tC[�>�1�=��u+�(pGΗ��s]R��ם���'yGZ����P	3�iR�H��t�!Eata5�����	IŘ!j����}UcܞڭM�S�&c�|\ԑ���4e��B��ޑ/Y��iZ��2Ry��i2C�����V�ds+����F���Ǻ�M����2� �&^��?�i�d�?�*���ծ13��lG��]�g�1<P;Xe2��`��x�mё>�j{E��.��dL�S+>6U����jP{�3 ��:� ��z�{�Q֘_yI@���(ބ��3Y��u�k���Ԋ��RAԖ��,&���k�4���~Nz� c�穘x�������Z-�qT�����Z�U�V�f��U�6��%��W�q�S�]�̷���ٝS0���o<Pc2a����C;���]Q.Xh�S��Ky�{{pI����d������e؉Or?u~�����w#�7��R�2��.�ٱ�R�
�ؖ�j@#��]"zw��HM�Y�T?oA�RSM �=��2@�Sͦ�#�H�F����(O�%�*P�͜'
[�����g,��3�SL�b��2)��������3<.1V'nd�4.�s5ChOq`/�3+冶���[߆�p��F(��)H�����q�?�v�͜')?(��dŬ��X�y2:�,���خ���9BX�\$[�)�Q����A���۴������P3�s��8��o�ܚp�>5X��3�����g�'VC�sd�������u�z���2KŁ���
�9���=a�ӱ��T��6Zq�)X��VЛ��C+0�p��C�e����u���vR��(:M
ʷZ�3ٺ����l������ø' ��v�zҘ��YU:F�P��
A���K�1o���A���&��*�8vzVeeLz϶4*榣�H^��L�ОRi�>p�祐�?���Y`#��$ؤ�0?)"� ���ݰlQv)5CS��*�O�˺�tb����:U���*9���9} ǍB�m)&�v�e�ֹN9p�2u	;ȱ�k�;�ye�燕��4�U������X������ �=d����?�B=�A�2�r{��v]Řq�=v����_z6㏣����_��ļc��Ӽ�M'�Shz���f�E#��o���P���4=C\����;�Q�Q7��"�eP:Z15F��Eڙм�������w;�K5m�UL"�A�l���v^�� R���-��g�j:n��fz�ziQ�0Ʌ�nC]�mb�@�c��=���;"��`���q&|}���si3�J�ZWG��m�-�^�����"|�
��VF5g_ $�Q��!&!�M~Z���P����DrqƦ��3�;�R.��L�6���B�Sui���
�M�BƸ�C���Ş�q|����D��X�`�}�DkU�_쩦��>3]i#_��P�A���Z�g�V)DԤm�t+L�h�)�7a6荽�`^~�fTf"@ͽ:,��Z�T��9�q!�չ�o]X�墨O��[�C�Pc��f^4V~��rd�F:��?Ӎu�e�dr}H��\�F��=����4�L ̓�(����`�N>s����P���	G��O���{�Kh�I�h�=���H�[�M&[��!��qj�T�%۩5�q�S1m�I������{������x[�*�	�F1��r����'�bq�R����![E"��Ǩ�ň�c�J�*���='4��
>��b]��l�>���Q+�t� e�:�{�G�W�����]���n�*AN,jL���kИ�Tm�F�FZ+�Ň� <��[/E+�H�p���~gʗvRZ�Ѹ ���dp����|���ݖ�-�U�e�B�/�9�Ŏ��Ī�!�hT�rͷ�ل3��_���-�7��~�j> ��.���l�y��πO���B���*�uG� �_v���9#0�! �����6h�d�'�{������
����;�3kB�N��اF&���Eh�9��r��{ξc�"�z�ɺ���2j��-�ZyS����-�W�����դl[qE�;��+�S ���k^�tyP5�3�\���1R����ٛ�����t�PJS�L��#�X��D�D7v۸U�1�$b��0��0�����G-�f��D{W/�����CN|���/ �X����U��7�}�����K ��e�����y-Q��C��#d`{۟z���!S\��	��K��h1c5[\�@���<3�� ��$�Cqe[�(Z�����z.%�mx���Ah4k����V��Ś_��Vr����d����Dic,%<��=�	�B%BBfxxi������4�ҥ~B�O�>aV�����F��m$�:�����:��;�Z�SI�FXL��S)�Y�M8V)��m���.�c
M@��PN���wtB7�-TD�u� ���eA��E`��e`�aBt`��ǭ����,��
�۬��	9�v��������S���c�D�#c0b���wxk��W�z���d��#�\/�D�O�̀qX����*��5�Q{+��@��F��%s��p��.��sV	�688�10�1��Ќ�UP����*朿"��I�U���V���J'1%������K�>z��L�'gLY%���'���\�ܢ<޿}n�a�m�<n��o�$�m_��z��-	�����{�WK.�ܮ��_��ٞS��{��g���Q';���U���~���]�\��y��n�ur��ޅ<C���\s�K果'|�2�a�Ç�m߻:N+���:"W��-�k��l�$#�B�r�nH�nD��`��>K\ ��~�Z��L;4���fxH�/�S���C�ߚ0���h��1#���g�oW΄R���a�cE n���0ǩ�j�"~�ܿ�螳�[�R4�'z��/�H�fT�-;a:[!��Ӳn�ҳ6�V��qTo����f���Z��˝�Ƹ���եM����S)i�\�H88�4��R����1���ʉס⭵zy(^�b��/�j�BG3xѿ�ձ���yT�ACTqJa$D�6޷�rQ�oQ�t)4<̳�b�"�Bֱ#��3O�#���٫y ���23�;q�Z���h�_�d�a&K�Sy.Z�oC�X�(.2!'��tq����x³���G�P��L�G���P��vS���D������sne��R��7�X,���I�i�Sf�䁞S��H&�m�����(+]�`O��Q��PdsK��1� ϩ���Y�y��~�N�(e`[�M�c�$�%J�exxx�8Y�z�ǆ�?�u!7��H�^�ӗ�s�����ԲuޖQ�*}u��j�
W���EMڨdU�TrD�29D㥈L�5?ړx���u�ҁ��:��,z�s�l�[�y~��OnN��^�(۔Qڽ�=�!�
�\�>����7'&�!"�9����!1�<����= T���!i���"o�^��L��b Ĵ
,�&�;T�K���.;%�"Y�&%�yq��(�<��=�[!��7]�z��q��Gjh��I��T|�"����I�ݕ�ć��Β�%[vZ#�E-��m4Pq��rW}��ߔu�=2�[�' |�|z͗"�ԐZ����K>�ø������5���n�W�CM����k͠��iռ�g�t\I+i]�)�Cw���u�$]\�W������-|�'���JL������,�b=L5Y�L�)�vZ�Ԕ�1�������[���-S���F�2�!�1%&[��D+�kP↞���F�52�H;�M��zU>l���#�Rw>w>�`�������P])����d�T�+r���bN�W�����38����Lv��-G���ixy���i�g7�i�IS����4>c��?��Q�C���r���;t(D�@QngL��9,��hk�(r{] ��-6C�c�jD!� ɯ;��z��z�R���m�m�BBT�һ_�,q�s�m�o`Vا�-�1��y>.F�0١���0~�s
��oM��8H��N.Z���M�o��!ݶ����`&�|�Gp��[D��bN� �酲�gIo�5�_�Ӄg�jD.fO��\t1o����o���T�(�68�H��Gk�lP�՞̸}}���eD�'��{�ub{p��̜��3�fme�1 �+�y>��)�7�|s0¯+�g]�|��>�?]Ѽh
e��&���b���؃�=���GH��tP���(���l�0�K��e3��G6��,�O T(S�ٖ�l`R�~5ֽx� ;�D�G��e��	nZF���@k��n�ne5�{��ˊj8�C�c�S�>j#>C�%ځ�O��F�g�Dg>ӲIт�F�9��R��Ŝ� H��3���K���u�w�2����h�hO�{���M���� �zsۄy_Ԃ�ޘ����,�Y����G��b���\�6F��R[��c>��Iff�]#��4�.b	`
�_O�;b���DXQ��ĉ�Z�D!C�8Q�
N���3����xټ�����5�Zվ�2M��ŧ�;߾��{����gߢ���y�R� �`�����
�R1aMb�z�o�?p�����3�=��ac#��[	��v�";�Xɝ���������RVjj�b�3��\���>5�� ܜ�uD۳I��*��g%���^�1?�d$���}w!𸧡;��U�jK-k�E�L�I��.N�5kM��j�bY�Ilؤ��X�1IЖ�NPJ�,88ɑQ�@�9n�:#�<6��,0x���Zb .4�rA̼�b�֯!�xԤ��_��n���%��o��}0oXߖC�+�j�ﷴ�T�9�_� {F�YN��\�L�Q}� ��b��zO
���v$[��
�iAL�I�0s�Y�!�E��xá~�!�r3SAg���9��P8���ې�!y�
�f�`u*|m!s�8�fo�����{O�d�g�l�h�U�࿲`��99���(�I��Z�w�'W��bY��)?G�n���Z�7<�u����r=ƑY�"��yu��D�K=;+l��[�._�j��F/�mV�{�*w�����YM�(=��F��o2��jZQ,��@�G,��/���[���0l �����J&5��t��E�܆��N��N�|�� ���s�3 Ҙ�v��m6�b���F������c�O��u�*�B��2����r5��ڵ�Թs#T ��Nq)E��j��
G�#q�tI�����f9e�"\�����O�m�\>3I= �~D1 o���e%�SzP�c� N�p㔒2�MsY#�<�#-@U�؉ڔ�5]�x��f
���n� Q~�/)������Vf�,�'߂����1�:�P�[m�����.~a8�A�M����<���/ۗ�����hc{���]Nr����U�����������0#����YUO��5��E�G��$|��JGq"k'�R�[����r�S�Z��1Sq�����r{��T$7���7M�q�=+���T�p�-s���f��G�L��[�,[!�f?��$P��v	շI�{���|)<�	X�nO��0�����GF����^�!��sRc�����鉣�T��{�k�JwN1���|VD������e\DzK%�e_ ����v`���@��]��c~U��n���؛�o��:���j~����	ͮcWT�a$��b��;�x6D@.ҭ�2�T#^bd�h���G��ȉza[��%�Ӹ[�j��l���s�}jn�k�#>ML�\��&	�;p4�%L�y-��|��U��[QXKOR�ka��БK���\�ж���c��������s-�t��0S�8��X���$�b���	G�x�%��mO#Q�3�ů�g]�&�|��G�y���R��[y"acJL���Ma2�]>!+�ί�Z}��'+�ЖO?yU�/�},�	��[��Y�f"�7��-&��[�W�(" *ڜod��������8\Q`���D�\�s��R�{�i�Ϥ"���������áH	nf�\��k�c�p(&c�ȁSO`&��_�)J�$�
����O�Cqn�J_..��e&�G ���	Pam��;
�� :(l���B�D8_6"�0W]����"�3����.i��Z;�=J�02����z�i�������$(w':���JY����}1�Xx�'pf@�MDS�h������.XҶQ�"�Ɍ��+Ng�1�ÃM�(=��ti���ƃ��.?�^�%��s�Β�8
\�*d|��6B&4L����0[���.�H4�g��֯et�u�BC�+L���(�ԣ��\ؿ����7�u��x�<��l��t��L �8�g�$k!����CW���m�_�zM����Ya�E���-Q����]��ߍf�sC5�K�?"����˂��ʱ;b�H���,�>Ϛs�O	��wV��Q�Z$!�{�f�YKH����y]��~��4lcn4�)�?X,��#�K��B@�-�֕gg�
��MӬ�HT��`�;�g�k��$��e㥲뙼���ե)��¿p :��zͮ�4U�5����,$�������?�c� �
'��V�����g�37mhýH��Pu�N��"~��K�k�`��^������YGzy�8��􌧇�i� �p�p��2�%å1f�7н�n�R�reW<���ĉ���u��q51���D�N�6i=��s*W'�#*��W�@��LJ�?�,�^�eT��Z�Χ�MM�f�D��[����K4�m��jAϓ��:$�G��ZO_p��{UA|(���$�AV��bj]��9�R���:HR�rX�F���R���"oznL�M\ȹ|���S��E�P��?[b熊$��#8��hXy�E�P���e</��*+k���:O�����U�{��7R<��P��
�"��w9�(����O+_]������)ja^8��P"�|��Q`7ʬ����LCd�]x�˽:���*̍ɕ$\q��m7c�+4�7�;�)�6�r�k��~�E+7�C���X�'CK�2a}6,���#	#ٮ\�72k��6|�=V�=���G1y0�/�2 �ge�T�*^.�t�V�������`����M�*B#͍$�eK'ʮ��f��gF�& ���3(��)~x�Llw��DF���`����p�"�"�e�:Sٝ(*?,��߀f�m�`.I��ٲ?�_Ж��Ӛ_���f"&<A�bȅ��/���ԇsO�85��뒩H.�?v�n��g�Ri����|�f����<�"D3�];]�|Ud"�����y$z�b�4��I�S�ʂ��Cڛ�Y俿;G���'y�U��F7�������?����Y��>nñZ��B�(횥b���X-9��6���x6��Mh�"lf�\�tp�B��m==�r�? �r�~Ę�#�X���Cv+�J��I5��dy&Y�27���5v 4�w`c���:�v���[.YG|�s�z/�Ԯn�7�NJP�M��ٶ��3N����2��[=ԲZX(>6�s����x�`t�QJ-6p��x�l "�e�4�Ә�޹�FKI@N�������}�!���闂�e��x����}�$�ē*y�FA�㿂�ǃ���]�{JD��J)n���x�o��k�a5�?%v��H�G�w��@� �,��LP3K4"���85W����Jy!���8h�z�q�\����e� ՜�`R�lꖹ�Bc��MSc����D�n�V��q�!�e$����"QN�'wQ�.��ɧ#Jxu<ES���X$xz�O]e�g�w��A]��:W�h�*8�Qg��� ]8��q����WD��o���98�X��8�����6)�����u#�N�w_��F I�O�q�R���,��"b;j��������{1���OR]<`���k�O���ۮ���������v�XU,����"��:�	�D���������+Y�Gؤ�H����"T�>��?�= x�XR�������j\���V�7��8��CWߏ���B[�zX����N�����57��sL6@�kW!1�N(�X �����30|;�.�(@�p��$�`%�C�`�<�3p�У8O��H4���H{o����N��vL㯠�DԘg�7�kW�9�������"�h����.�Ѐ�8m],��؀&A��t�����5~f��m��? ���	R��������E�;M��4����k�J�:#1f��V��~��2���a)�s�L	��r�=t�ށy=RP�Q�P��8�<n]B��"�f�Z��B��� H	ӥ��������F���6����+q��l1��V�W���(��cZ���E%�s�ց."创�­I�*Cy썟�2��۩^c��UO$^-4o͟�!������a����[㕧1'�%m�G���6��ܔ����K�F���RU����MFE�:���<\e ��Ddq�^[�F�yko{�&�%�Q=&VL~&=:.����8?���P^^21�l��=Q�B��6ɛ�a��O������4W֌�Zl,&��"B�g�k���0��@��?q�A~F���JN������u��]�1G*GWU�b&I�&�GD�W�� ���=�tk���/&�
�椈�w}9;}ṡ*c�U���u5C���^��gM]4�2�[Q����eV�mA��W�nR�F?�n�~q |�E�~�>�4�
�p��d�j����MTU����k� B>�O^:ѕ@׉2�þ�:3�e�ۓ:C��F6���22}�ѣ�v8��oHP��r�d�o�a��*��/�����O]�_�Bܦ�fAӀ�;��詺��]�|Ss����h�Ś�H8�b�x�b���b=���m��z^���[[Ѣ�`���IS2�h����I\ƘP ��|.�����$*ȑ�Y�]@��{,0�1��%����Թ����(�Y�O��&iy�?����Y�FU%��rF�� �U�M'o�%��MyLo�$��"��,n?n���h	p��s�Ns���͋�l .""ʔ-���N�>-G%}[���nʺ�"��o�mE����y:��5%��L�������6��>TEՉL��m��Ze"W�_�O1�)ݎ>@vy�lgU����t�%�G���l �ll�$`�^�%�@�����+�P�f���U���ߪ˨=e�d�W�" V���A��k�$^T�|�b6
�#
�SG?΋����f��#�����Kұ���,\�Z��2Sߢ)����1��?ô�&��q�����BG$�R}5 �xp(��I����o�[�0�[�&A�	^���P�5�Z1r4��P�����y%(��7��1*��{V�%;��T����ʖ�1%2:�J	� ��Ȟ&�E`Ms�/�]�'���?>֨����z���1�d�yL���Ϟ�g������. ;���C��~���uո
.�I�L��^�M	:cCԴ]~�4�o��� ����V�E���&���$�޾W�+��+H�O9���~�q���߻sOÞ}��'D��'�G�Oh�e%Ti���%}W,=�)dv�hR/���/�)6���5oks��$�ޙ���'4ry��!�$��l#�Q�J�E)��#T4Pw�@F�V�y�����-յ��Ğ�_���V�����R|������l��ؘ�(Ov�6���鲄4�NE^���S����g�u�]	LP�Z.���vg�����
���N�,����wg-}ż�3{�h�~T�ܷ�ƱrD�.���r@���dW��q�R�*��ʁ �k��#)qs�`�E�L>U5y�ᨖ|��|b�����V�F�<�X��z�A�F�y^�C���5J7{yba<	<dዮ�i?[ۮ���P	�D*1K]���H(+e\\j�h�{���T8\9�?,����j;tK�m��6�b�M�������$aâ�uwC�?JWΊ���=����<��ȘI���Q�����K�L!!�(��;��wQ�A
L�t�WX��ʓ��?Hg+	�-w��
�u����K%X�{B��3�c/���E��D��˗}g��4��v\����EZ0ٞ�`���w��=O!�����I�!c�mAk�^L������rwjf��d@m�Xc`iVM1�S�
�|���g��Z�Z���� ��%� ���X�UH@��P���Xnɳ$��>k�Z�Os��9��u#[�*�l����D����- ���[p��ll��m�s8>�ԿP�a�> ����J��/��}��h�7���cq��!�P
G]��<Xr�~�������58�k�茸��1���<v>�b��.���s�#�c���b��y�f,��L� o�W��!��.\o��	7�j�r2,�6v����˻ "�2��zU�W��U�d���-Ĳ�]| o�3q1�M��fpK�,��dz����%``&�Q�&��i���`5w���_ �������s-��(����pWH�"�ͺL�[�֪���A��޻hj�i����X\���>��Veb��1��ִH&��Z�ﴈ��C�v���Mu�e��P�hL6�� p��]Xt]_WO�i�J;2m�4N�˷pFx����3�K*T�R72yk�-���y��e�������s;e���Fc�Ql���b��|����Y��K�~����)
�	Q
��L.�%g���=��bVs����s�5ԅ7l�u	��H�0:T�qoﶰ{Lm��,|0�����������HTDk��#���ykX��+S�7�u�L�>���;�L�_�3��0�qG+1���_�8q;�o�g)Զ`�p;�B�ߞ-ɦ�����ݥ�P����W@v��ipŁ�ژ�E	����P�H���M�ۤ��b��BG�Q�h-����-9V.������Ǎu8**�o����Q�%gR���޺͓>�,����Z��ί����Ie�Gw<P��&�T��D��>�C�Tdf�Y�D��aT�@]�a�o(k�~l ����6p�2�r{%7��d+�Xٜ��Ť���J�Hƿl�Up���kUv�(��5�Ӣї"����+�k�'�%�U��9�J�F�2��ژ�<륿쑺�w���g#GFUK��Q�RIH��Pg3»���׫7YR�V�p	C��q���я��v����۳��d�J`R�[M�"�>'0�K�=���"�~���x@���&\�BlFp�lK2�J�+�����L��
�\"���2C���/��9�ى�Gu��o�K��J�����X.�o�PG�Z��>��yJ�!��&D��p/��if=ʉ�;�%��Htq-g���FW���Bу�hO*<��IAtT���$=,��Jz!���^�x����C�ڣ�D\������88���|B�_-�u?����~ݢ���"��k��:��-#�:��Li�z�I:TG�WDNY�� I�C��A�t-9�1�Q��d�m�MX7w��?�����V�F]籤�TY54s5�T��vn��,����Y��#���Q�!ni�M�nڪ&J"���/	X2y�~�1�Z"M;l�@�7��,_�";��9/5@���ѹB ��Id@)�:��!�J�/|>�K�A�Cÿ�W���E�,KN�	9�����W�����3�T��N�'X
��t�g�N�9<~�k�V5n��n�p����h��� �{�+A��^�G�5�_�m���|��+N1�Oa��\:@zd"�OpN�Ņʰ�Bp�~�� �Ӹ��SMn�ޮ.U7�T:��8��g]n$.PF�a�����*D�K˖J�E}aD��J��#��^1H!>�U�`�]yr% �vm�0��Z��*�A%�t�X�f6,h�k$��g�ď
��O�3��߾���A���\�^w:N?F��ۅ�;eM�V����
����}x��l^�������̤�I.+dˆ7S�����y��߭���K3�8�V�Oc8���`P1�[
�_[{53wӟ��@��$��#f�:_��;�ď�.]�����N�S��@�V�k�} D�q��)I1�����h��0�1%yxh��o�
�.3��� #�c��loƓ>���$��6��נ��&���idΏ�-@����-�y4W|��R ��@U����������$�X4�Ϥ�	L�!��*k�P�a7���|�L7^ڋ�޼:	��҂�1+�3H���S�d�3U��Γ8��62{cEͽ�>��[�S�'�?�2�dӬEu��3/�OM���Mt��Q<5�)��Q0ە����*�����i>�?	�=���;��zu=��.�9�;ObF������<)��vc������ص���c�_t��`r۫���X,�����Dq�-w�:ۘ��c�]m���+X�o�yN����ԉI��R�A�w)�x��S�o�BwA����-��/�Kk�� rS ��ͮ�w&�J�� ����d0$;��_�T2f<�U�X�\���HqIf�?�;aP^#�C���{ioT$�.\&�{�L��߮�����jƜ�-b�2�k�h�y0	������jO��$8V�O��0D�~�v���ȵ��^�}���΍P���ĕݫ?�)��Z�U�9e��Fy���L��.��&9\�w�k6q5E�4n�[�K6ѵf��
5�w�� �)�jY���<�'������ES3=��u�v|a�3`���%�49���0.�@�]K��|�[#[�RaX�8w�MuD��.`�[�x��.�u���ֻ�;�E|��P��?xG�u��\X�V���s�S�����4K���(�����s�^ӿ���E��H�S�=���$��;��n�h�����<h;?n)�2W��3JkT
l��V�mB9���KЎ�MmH�����ۓj�A����H0��ØS�}���>�ô�r��X�}3�¡)0x��'��mtt���UHRBm"��<I��~��|�cWAe��wZC��Fc�Gں�c�54c��bO�;��o����C�-�p����3����'�2�L�ZlŎ�Ykj&{�j:H������c�oE���;I{x��������`:ʍ�XJ~�DA��Đg��-ΨPQ�V��6�����i���h*�u�F�.�A��rAy�_��(�$�)��W�c�&�i:�1�/f2�=�4��-�V��{r\HN־� �#+��2�#��C�S�N>��bE�8����s�"�P�=��iba�p�SB°q�Ȗ5�.��������8ǅ:����^��z�ѐ�C%�q14�kS='�ҋ,�e=�e!��="R^*\�ܸ�E5r]o�/i��m�ʤaDX��Zσ�;ܽ�#�6C� n��j����q8��;�-fqa1�amn+Y�!�|k����m���z],�p� E��=sV�����}
ӬX}U�kD/��̹^�FU�Ǟj�AzFS�h ��C�
�$�U"d(�>��$Ӈ�*�t53��bI��꼸Zu�9�G�<*C���as�63�ٺD	�"������'7$�+,�I��m��F���x#r���z^W��qƓp�W���ͦ�4�p�7�U��v�\���䋙�&C�4��D��p� %v�YHB�ml4��>��ҕ/�5��bR���б�"Y-x[���k�M��P�z����dsNC� �AG��$>��}��� ����8].s��?28��8���$l[[
�Y��=�[MmX�� �J�#j�?�om�~4�%�RA4��g�	<��1C^7���MY�������QH�:��f�Vƌj��ې�\����A���P��ғ�؂I�
�w@(�z�����ܧ�F��?�QQ�e~�֪c�K��o�Zy.�R���f?Hʲ
N�W��?�ﰱ'��7k��ǔ���%�{���bQ�WHO����
g���=I@����$������K��ؚ$�Uv�1@_RA�����/������p�44{���p|6a��m?P䮕���z��xИ�����ԕ��R.��3VM~�i����H06�q�<��K��]a��bAl[�Ȏ��;�i�+/a�[S�PW�"�F��r7�q��:�b?�)ީe�{�\eU�rD�B���3�1��ܳB�m�J#L��`��RWa��"O)���e��G�#�'�b!G(�6�����l�f���M���Qf��s2�Dr�y�=�����?�e�iq�M��k�3;���|3~�j����h��Ab��}cj9��.7"�|���Z��R��ӽ����9����<�'Ay��������>h�O�l�N�I����l��=�O��޷l�t�tX{F�)�t(�n�<@��7�澻7=�W%U�2/?�q8K W�$cÄ]@��$�%�kA�+��+a[�B�T������4+����
�},1ia�XA
�"$���*�����Q�\�ZJe7������Aht�ӡ�m���k�#�퓀�Wh05�YB��U[
 _�s��X����qQ��(:��=�����r.�B��X
Ȫ��{Jz�mN֚2|���l��>�4K�m�-��4�*�)ڻ��ڦ��Td�%�t>��z��k9� �6AM�ݎ���{�q���e�Ft��5}��LSV�o
�|�x�R�~�q��aUA�v��H�q���B�SL0X*��?���Y�e[���K�Q
�iq�JG�oP��˟J5��y-�AX��ψ%����L�ڈ�$aϳM^je&ۥr�P��N�*�mMEu�#d.���Ke�n�{t#���2�f nT�Q<�qd�Rb��
����j����'���ྜྷ%b�v^�9�q�b=d�r����FB(��G�t�8����_�K�na�$����ʗ�^Y�>)��	����s����u~ۀ��C$�x���͝�������E47Q���qR(�/)�b���S�B�z|U(e]�C03X�&u?�O#�7��k+|�;q�U�����\��_�=9�ِ����Tȅe�ߨsk9�Y�Vy��
��FU5�e��;���d�/�d�u5l2�|e�v�m
�2��h�dsX�8pB~!�1-ܟ2�v�y�H�.0�����㏽@�^����C��p�/�6x�%���rd�/$]]
Hr��].:�	�P<�Q<�~��DE"Eu�gd�o�4��Fp�_"�k�:|q>�7[�6{��W!';���d�4���Պ�I�
�:��Sh�Ӣ�4���s���.A;�d�k?��@mTz�?�G�C����s�i]��T ǁ�U�r:�s��.�^��1'�{��z�S�"8�H�k��9�\6xe1� m�)p��lGx�1L�82�)$�cp�x���rd�;���F%(9ˏ��*؊����z�ҤA�����~�pZ(�8��N�P @ .�������!�)�����F�0m�?4��*��ZGC��:�1`oD�O�)�3�Uk�kN��<(v0i�Rj�ՙ �Cs�flƵ��9Q�����B�0J�w�\&�
��E�'	���q��9щ�#����R=Y\<��Lf��}�AH��k�p��:���搢�>EPZ}0��U�eѧM��{Y���nu��o;�'�9!֔?)~��1ֿr$^wer�=�9���0Ų�+ .K��9Bi��Κ�X\�q�?(�m�F���Z~�]_?]�M�.�	T^\���"��@M�Z�R�z��(�{d��cީOc�J��V�O'�<&��6P���lI# ���X�����,��ԭ�O9�����kb�Dd��g��9.l���ŕx�c�V�ʞ��|\Xf��pL�P�,����ndZ�p��%�u���ȉ{ou�K�ܿ̀��AիBԨ�ׯ{���]��c��H�OF�����w޻��a��~�,�ￔ�VLvǇ� F,�B<����<����[��'0�W v�֐�=C��Uj̷�t��F�:}{F�qÂ��9��f� �!�^\"^'��
o�,t�7��{��JEK�����	�`��7�X����p�,gn�k��bl�m���1+�Ϊ����e�DQc� �Q`o��&�@^��Dl�e5�Zju�q�o���w��իVM��A0�m\_����(�,�u��^�'�J��P����C|�"z&��ډ�?GS8�S�;f��2J�p���<Y�4���� ����l-��rdR���
�|���Ƶ���4��D��"A����X� &n����39�sz�*d����'�t�J݃	�w`M�V��@ ې��.V��XMsaR�q�nƨ���.o�U��b�{���
f#h��{�	�ǃ`�"����<C�g�ւT��s����Xa��J���]�8��
��Q�.iGI�m�6��l�o/��'M�x��	�w-�I� ko?�DI��|��m�Apd0C$���l驳�J�O8�p�LCw��}	d�Y<Q��ĶΟ?��HX�<r��Q��r�j����=%�+���TC���V���J��t!��Z`ඃ2V([]��Aٟ�Z�;�i��.��9*tM�Q7�'�ч��n�&�i�zv����n�3��q�{�*h����Q��+���B��౿�/L,�a���
bG�������7���Q�sXO��xN��o��Ӟ�s3	KB J��.�Q7[K-W+�3?�:�n���9 ��<�g{YX��4k2�0F_�Y�+��w���;�v��%�����#Bn��jy���.NFI!-�x׬���Nz��pa��p��Х��Jl���m��W�H���~S��M����shx(��N��w|ӂ�U3�)��I��k\$P�vu9C��K� P��VL�I&�1׵$;�ݦ ��L��}��A�#��?Rަ�%�Ju��"�3�)�!RJ����_sze&�e��t��5f�jFR��s����;�,.�Ά�a�i�>ў���U��a�+\i2�f���y�FB�(��g�pR���5�1�èF,Y��'�Cg%p4k>�#ӛ�k��⛗P[��� �P��ͬcI�fp�l\@�ԇs������s^%�.�2�ͥ�<���%')�&�XΒ�3��$�e4�`�(��|н$�>�?ǼY��#]WtL]�����nK2����#�	AY]A��Wɖ%���d�֧P#o� �ˍ�GSGz��=$�,�c��pJ}�
���{3�-_Ɲ�>Ȃ�N�cX��}���Ta�O���A����QW_Vf&y�e%"<Otk͙��PЃ,���):�a��Gk,�Q?H��]R7��S ��$"Jx�,$�Q����"�]��S�i�?
ɟ�N�>�hI�����"��P���~���x�`�Lಋ�Pc�W�L?�^�X5WP'5<5�V�7������7� �dZ?�)��t(-j�q��G2؄x�Jof���~�P�tr�kɾ�=�Y�G���%7�IJ�[�9�P(g�	i5Q����������W�w[vx��ف�g!QAƄň�CB����զ�^)�~_4�r3��-�K�������W�&�C6��q4���&A����a	�@D��j���j#�0��~
����0!����]�q*�C]�׬�0�9J���V�\�*�5��t}i�F'��L'N��SWJBK�;(�u�S���W~'@��ث�J ڐad�7�*�,B#�Y�;>s����Ez� ���'��s0v�>&������t1.���J��(�_k��L����7�rE-g��6H'9�;���I�BJ�3ȫ$5"�K�N��I�����_*��4�9og��QK�[9�M�T��PW1�4�6�CC"��R�2#6')^�2�p.���(t��|*���rO`�#?�ߤ�2G9'��Ѡ ��H������oJ�F�d��nj=IK��4h֔�V3��O������<2��\��&����:~�u+��<�v3�+��e/y^[~fQ=�3]�������2�$t'�^k��cD�+��l����X�z���R�22�KG �n��������x�.R8!K�����3���$��j˴}D���\ �6���{��d�p�N�O��3�N�CF���?�?��4�\]*X���,�n��0Ha��D�9�C 9�q��?,{Qll(E}rd�����>$z�h�rV������2�B�lj�p�fFV"��������JS8����Zl�_�� :�cȱV�y��n]��P(ա�m��K [���` >�2,^lͤ����t���M��=���t�y'�g�Ii�)��JE�����́F��Ҭ������v}��c@�lIF�����5Ց���)fu��!D�7#���ό7|h$�Z���;�!���1�5�ԯ�O�3�
	r�\@�_+t�JP�.�c�$�д���bɹJ<�����J8���DO#���p2jUv���Rߧ��m�ͤ���ӵ~y���v�@�����Ț�Q#\oy�z��E�䭡�c獸g��~��K>�C��ͱ 3���{�3�Pz�>eY]")A�5��mQ�����%	��%�3���j0�l��\go�(8]T| ��=���oi�g����A�"�m��'!r�+t�����=O�H�=��1#q���u��_� j�CZ�!9%�Z��5z�*ڭ����|fM�5��{�� Ó;�Z��@��i�w����<���g�
��$k��,ꃰR���4��k�f���[����\���jD�2��~" ��zi�P�r#7�(���-�i�^�.S .-H�����=�n����KaL��9�O���ͥN�z�HO91�X)ฑtJ<@$���;�|o���n˵Z��_�p/ ��*pg�(@=�&���s��������**���3�u����̰&�K�E���f��`�Ω�������9��!X`:�c;�R=G�Mjc��p	��A�+��pDqC:3�@!�Q�Lٻ_�h��9�.�`�4 ����P���\�"�>�!ѕi�/ZCB!�U5Vp�1�/���x[�ͫJ�輋z��#�A�$5fb�\'	DOu3���o�kW������̒4G͸�Y�w��rh��~��Ʋ�g��$ڽG�j��y�H6I��GK��|+��gUj"�$VRv���3��S�_�A����߶D<C`cR��N�OH%EP�'�ɔN�;��$C�n�w�zB��Ĳ�]�y.���J'�!�)�W��S���I��gm��諙�fa� ��diV��`�-H�B'N�e��Y�GQ��u�����r'��oJ��M~F�r&�w�q�m����1~͎?��Q,vρ�6�z�rL�:�:��y�W�;⊱��3�|2��G���#��~j���&V�-�T.�f4��Xh�ƕ"�"�H��mPg�%KU΍��QdKR���:٬���̘�KJъ��d)�D/��ƗU���8����c;�X\�YNG����>q��_���ߐ�×��2�F�׭L7�#�P�b����D����/�E�R�=���sK��=�� 9��Hǡ��4^�R p7%c�9ʣ�S�����Ú�p�l�����LQ2h��jy~�C�b\�>)�^�v����@�=�iʣ��㔲hѴP)�^��#a��n�,���:���tV��T�D�P�6eB��
W6�� j>ڙ�.?�����(�c�v��=� ��9� ��� j~�K�e_�Wm ��cA��Ჳ� d��]^�9EE1y��j	�٦6ѿ}];�I��<�K�`n����յ�_����Ӊ���5�y(U<�u�c�k��O_sK�yaHkÓ�
�:�=�a)/��nRB��jSm�P�xT����?j������dc�s���e�0�""�H<���w�u���wHS,Ug~��\�����t;�H��p�ߵ݋�:Sص��H�j [�j�u~�Z�^	�.��J@/=��9)�M
���~�%�[���
�w(�6�N��Dxڹ�kR����vۦVj��+\�?�Up��+���3�3�(�+eql+��3<f��-L�N�x��c���%�_K�y�T�0	���j���n�
hq7i�S��~g��t��#�A�L�A�SZ"sj�r��s�']��_��������`��{�6��'
��Pj�ܹ���͈��§du�P��y�I1�C,��a�u�s��R��<���[[��y��IF���k��4�gba�+A���å��Q�Wr��Lm�95:�p��/_'�1A4�m����CV���fY��\�9���t'Z�@o�<ETO�;_�'��Sl�4��D���d��9~k��1ŕ�<����lnO:F��!����"����2@�X��GYf8n8-z5�Wps�3�A�1���/D���B(y��1xPi� �\t�b���a��ۓ#��k�.=K�-Bz�{\(|��"b��H $Em�I��"��L�����q�U �~�OjFң����{Z?����|#��au���`�k{���9����.7A�����+_�7'�\>��brB�;.�S�dg�z���R���Џ$d�@���A���ظ���G�z�ڟ�[8��D>Ƨ�X	�
� ��y~q��I62�hW������*�+F��z�%�4��X Z`����+����i�y���wf�7��0�>yl'�}ŘƉ,�zOlR�B�˂�1�B���0gŢH�ۆ=?�΃E����]�/V�H�<��㋺T��ҽr�J���tO�!���F#�q's3w���)�ާ2�8Ʈ�Xד)<�ϰi�e����V!���5v�
6 �OM�9���_vD�*�bRl����G�8hep���w`X�-��`Pl�g��}�wE����Gję�����fEw䲺>����d��
*g���?�N�,��%�$/���؆��n��I8�3�r���˱zw�&d�+)�g�o���G��M�s��a��5w"k�*�ٞ4D�g�����:K-�,�2���\Y�#��T�0�x)��ю�-�"ՁuG��2��9[���]w`4�B�c�m�v��j K�u�'�A�尷�W���+�9X����@|�S�5�lA�ۊ-K�	���%������������ʶOo���.�I���
�1AM�K�J�c_�q"�����?i�Y� [C�l�KV��o�cp [:�D��3���g�|�v��~�/���y��g���U�鞧w��i�X�.Β(�B�D�hq8l��V����0�ʬ�fF$.��tG�\H��ףO���+��<�:��K�5iI�f�D��\j�Xye�������1�#Y���>�	��眣u]������-i$�)��RfӃe�<�ғ�������BWG$�߇��[���CY?x���>��)Ą|���1��mF8;ƿ�o>w5���i���\�3�©�%��:��B-'�b���/�>��18��]� ή�v����7.<�d(Z����� z8�b�	T<�&���D��b����[��k���<�"-��uDOZ\:<u���������̺��G-.%6�W�7��G�!���{R	S���|x�;��/�J���H�p���$�f$���q~.�Bd��ǝe�h�i8۽ؽh׼�<aRN�(nB�PR�m2ҍ�.�i}(;c�g��X�}��T�W��&�^��Q�C�6��v�k0>c�ξ�E�B<L��&Ko �,T��GQ�x�aO�sa
ϔ�G~��A���3�B9sz��}�a��w�	��3���J3l��,3�F[F�8xur! �婵�E=<��ŎK��`W�l��<J��EI��������Y�@^�� 0;���Y�n���Y��8��KA�
�������he��.�G!�p��!�w�OS�c�z�5��D���syP֒゗�JoS Ӎn��)��+2X)��`�����&c(S�n�Y�?,g ^;p7�����1�N��h�u�U(���NI[p�?�bu��kFq��% �mӅkG��}r�a���/d���x`zy�b;�5咳e^?���i�/TR��h �~i��}{�u:0.�T}S%GAHc�[����'C��J8΅�����R�y�4�3}q�[S�S	�:Q�(M���"N�^_�F�����ʽ�zÜ�z��IzRg$F�Fڊ��
��&����}��b�Hi�W���Ȳ�Ck,Q*8�y���N�	PA8�	���_{���'�TXO�&�\��^V;�elAW�	q�'�x'SfzEŀ����!��cȤ꒯|��Ⱦ���Q�8{��%jMLb��V̬wx�������4��e&�U�p��S�����;&0�F���X&F"��_Z�Zr��
�5s�Cǣ�9��qˋ���瞐Ђy��[�63�e��Ӹ�G��2���3,-�ղ(钞��,��w�+�
�����5��~M{��b�:����To�Ew�"� K�'�D"9�ۧ�Co�C�������s�ŋ�Q�=��is�{[�MfǑ=����<^m[4��lmv-1\���U��Y��F��ZA���s@���\G����wA��
�:\����l*�E��/�i��,~"���H�e�Oe���7���BΥdw�SY��j*�~�udV��ct��pvZ���}�Ȉ��i����x66��z%^���@L"���_q.�x�fo�AYZd||��������iB!�[�K����u)������Zo�c�nQG�{d�n�c��a*<%`�O{���.��?V�e��YB�X>auM�&[�T��L���5�WR�F�,b�s�c(�j��Ohz(5B<�D�b�r�	��$�W�/���ͺx�������p� ����yC��t^L�������6�
o|��7 z������<0�Y��-��>��8�)��c���м�WU�/�%+���>�� ȵ����h^/�L榁�Wtg3^dُ&�y��2���QVja����}Ӹ�ȹa�^��3ܕ�::z|�v�8�Qy�z�?��T��w����4�-2|��ʞ�<�aB��j.�h�8����j��At���o��n�$�1ؙ߉o:K�KP�����3�W�}�Á�	���p�/�~��O����|�2}�v�ѣK�����R�ҍ6�����a�t�2�u7�7Z6Ilֻ��Q�������F��t&k�X��
N@��O*v�~�OZV���tƨ��d�{����Us�YN�������O߆���O(��\�s����(Q��2>f��1?�
@~��H��b�����j�n�m+�w8����~;���(�J\�ʣڎş�Z�`E��)��hP�yN�j������C�uɛ6x�p��T2��/������r��Ȅʡm����@"t�eaVY�/S2�N���ӑ8��@*>�n�Ƥ
H�a��}���D,�jD� 7r��U2~J�z��PN��>B��6uu7�M��_dg��M,��R��m���(�T��}��S����&$��~���@�HFz��t���V�K����1�`�i��H^� �d?���*ˬ���К�SX\v>"��5:����G}��U�i��V��u�)c�$�lo���&J��u0�ʍ��k�6<Skm���
�7W�{�Bp����� �U�3?I�Z\�Թƪ�1��ͦ'~�-QW��,��A��9F�:���v/N)h���Ͷ,��)�~��5:P�?=����^B�".
׸��L�d�\'����7�j.���}���W�Go�%�tH��-+v3���ű���~��ش�R$��.X��uo�u�J�1��ط�s>�z��g�����$oSB���<��A%D�\_]��k+����`���[�G���6Rq	s��b�D��,�x6��j'
}�f�>�[+��;d,p��W�Ɉ��Kc��9��X��X��@Z�,F��� �������g��qC�z!�HJ��.�����=�z�����^xQÛ�B��FxO��:�[f�&�K�P&���m|K'F��8�H/¤��r�@��.c�y%�3���K�[�s)q.?�c��[����|�ӥ*R���@�-2\6�Z�!.�[2U[V��y_or�N}�7�����Yw&��o�i��w34d^N�)�#2���X|�k5q�vsܺ�9��l���I��&X�nU[�Ѭ��2��	��3{���;=�{��.GP�'
����R"}i�O3������V��m��� �b ��^��O��|oE�j��k��
@O�<�cj�p�@�(23V�P�����&����؏iY�?�. �d�I��9�e�Ϗ��-aqO�\�$6�DI$���gj�����%ߴm�o��Eޱ��'���%4�t�Z���Ys��`�N�W����k�S�[��99x���=+��W��<ӊw9��R���z"dˀ.m`O$����0.���W��1p��G�j��M�> ':���q4�(�|N��EW�U��"P��oB4�L](p��oh_>����R���k�'"�4v���^��љ�F-�(���ը�U�k�'����z�p�a�&��^�9�ڻ&���]L_P�����P{@~��V\5��ʭ�)�9���z~o��s�q5�����[޼`'�ڪD��Q����k�Lkn��9ɓv'�����f
��}J��ol��;��t���i�φ�/:Z��ĊU�(߇������3�D {M�҄��E;�o���l��Lb��������%bw�~�N]�ʸ�'ZdR웊g�Cӝhg�B�F��z��
9��m���旤L�c���$6�� ��bE�;bzm��N��'�7�;�`zڝ����!{���U[$�.:@e��H����m��0
p���B����~n��,�\���������;�;(+�b���������`D1��y�EB�9��s�-���36�h��Ҹ9I�0<o>��slFH.�>����&���l�/��2NЕ�͖I\*�3�M�u����5'ĘnQ��1$>�0�Jn&�p��ޞZ� =���W�B��X��~R�=�]�)���BDᖳj:�mⷙ��ZM��,��Q؈�{0�MM�8U�ɹ���ڢ�3��h��I��-����:��S��}:�g:M�v��f���YG_ #Y���CR�-
��z��wН�>��|�W�#u}����~�� ?N�)8�b0D��W��ޕRh�� �v�lfm?�س 3	�n;����v6��ZZ��-Q�iW�2mU����5�+ ����ui��������S�`U��tZu�fᰡ19����x��9LL��}�N�a��D�~�u�9=��.�xEh�^�Q)P
@��zƓ��ج����j^��F1�e�N	4<����`7A��`�O6b��{�L�H�뾿�6)���6�9w��4h�C���]D3R|��GŰ=y,x�h!M�t�z�.�/�U�R���>�G�L��Y[%qt����ɭ�v�Nȭ�D<�vF!�e�W�N�\θjO�o�0Fؿ�;p�e�G؂�m 7y�� �`���������}�഻7��ڳ��4�y���A[�\ ,Q�7�#7�
����h�s�8��X���s�H�wr��X�8BiwV��3x��R3��c�!���¼0��j�~�d���?t�U)���"��,���?D&��Li�����!O8��A#��	�_�^$لl]p��D,��W�]8#j5�v�$i��M~<���2�����άD� �礽'���Qq�e�;Q�N���\�p�.�����l�>��NQ0HH{�:vU>���N )�M���B!?�Tݴ��Nw�d	��p��'�c�[ds��vG���7@^/�C�`��kh�4����pLo�ܱ�}�;1�}�T����[��	T՞�\y����� @�����j���%VS4Вe/�o��x#H�1P�t����J��FWx	>Gܔ:�M<���N{��s~C=	�C������?a���M��=yE��J�8��8uZO:3�����>�)�:qC$�3mc��w�ϻE�#a#��U����+���M	���m�$��;�5Ji.�#V^[`�e��� �L�}r�砕֫�SZ��sX�x^f���0�Ueq%�I����T�25��B�S����Bw�|x�C�H���]x;���=R3������mD,���4u��%�|+����1���:k�&�Z8d�eG j��86����̞���]���aUgq�O�l��5`>���N�[wEh�
�*�_�Xe����:��4���L7~�^ͼ-�%d��B�ۆJ�x޻��~�.3#�K�*�������0cЭ��vd�kL�N�||�UDf��Cw��#�Tq�aae��MJ�=P�E/:��)bb������4\uG�cG�:�B�1���~��1qhU�,�·�	&ca�܍|�"��B������}�Ȝ�V6P/���7?C�G��Ece]�3*��B���x#�آDM�߆=M���+a�g��{2;���~o��� B�� �u�C�'�+�������P4�������4\=�>�!W�.ZCCo/��J�"&�o�����.�h2j�%F�j��x��6s>�����s0��W�/�M}�Ä�?�X��+1���}Hl+�Z��j��s��Ltj4<�aU��T�ǖ��V�W��#�|Ąn;r?:�l�>��� ��y}��O�����Z�:O4�#�:Hױ�Q��M��������I{r�MU��fz� K�X����I�G���o���|]���79���u��)�i����k_Bd�Z�եm<�51�g9���|��js��aB
Y�Ǵ�Чk��ى�}Ldh_�LcJ����^���8@Nu�vw�6�6@H�H��#�;Za
'�>#zN1� z*�i���ym��
��aU�cU��=B�y�~��f�O2U{n�LG�W�Sw:��ե#ݰ��Ft��dNpii$)E�H��n�GoF�m�Ѯ��i�R�62�P����
�:�N��c:.�i�ǶڣEd�����%�~g i���#+�z}��r�������}!�zP��3T�3���9�U4�1Q޾��i�v�2�>�/�׻z6�q6����q~�H	?�C��<���X�YvI��W�&�[��vZ���g�^�\sv2�o'���p�K��x�9P'�0���՗R�$��u��@�U]����Q�p��u�w�wXz]3��'/b`�T�k�PX�Z��t�"��SP@�?+>���|/ۧ�¨�BP��C� ��1�����M!K��b���1w��t�ݣ�0���o � �@�hb��N���(^��w/�����U��{����3�)%���T'��4-'Ԭ�uq����� V��m��ġi�m߉�<H����X4�rªR������יn�v�Rq�ء?F���Qֶ_>�dG-�@�Z������`���v�� ����.n$'��0N5�Y+~!s?7Ou37j�� ~]U1�Ζ���o���=�O;�Պs��qUz�,`u~�ygw�ҏ��]jO�g�,-��fM���'�O��-�<y�;rG;P�%rM�9�l��ݳ���1���u���������:�=fU�￿���;E X�����ܼ. �u�ECxV+��7��U+
}W"���y3��3ڂ`|�fs���_�$���عl�E@Ӷ�;^�\̨������(&���W���!�
ʁ�F�=R�(\���ߊ�-�ܔH�hP������ ��5֜u�VA� 5��KM�DД�L����%Bj_ĨE�1��Zsg9��87��m�h��?�Ã~�+�E�^���/�Zvwwlx��c���+����D��l1w[�-� f~K��Y9g_��Y�;�O��1҃<m\���qM��O����R��噻z>M~�C6ՃnV�w$��6>~�Zan:�����̀=l縼�nU
"� ga��_�+�u6WT�-h������m
9
4�5ka���4�3�44�g!G�D��ҚZBl�K�
t��̙4l��V�������2be:�c�Sqĳ%��������埡ݛ�,^$�q���P�����MĿ�`#���5��D[��]uDq]���b��=�5B�+�������J~�앲)C��+��^I���y,��t��FBo���./	��,��!�o�.)(K�g��I�*�b�O&�-�����|�I3�)�pn�?~j��/y�ZYE�b����:��m����E�q�M�l`1&%\��R��`��-�̶Q�LM�d�z�cd,1X��^����VK�w�S��4�p���Rpp����zp�w%QT򧅒t궚X�H<�6�1�_!�y���t
u��^��f	��;e8�@T�z3�`S!W+��y3z9���I���n�|���v;�����f2:'�{2L3��+���&��z�׌:B�G��R�a�xQ���zG�J(�����<LgEd�ެ�0�9a<jQ[R�Q4W�)�%7$�yB��� �T>s=��g8g�_�w�ر�N�C�y��.A�[�W����)u"��)"��t�?=ڔ�Eޛ#F�r@�|�܄e�Y���n!��o��7�c5W\�� ?CrG�t�e��0�Y����1��)�*��go ���.u=����B�Xşr"	�~%a�զ�Rh�73���Y�"6�3��@���"����ҽt�C|���IƪWU�� {��5G򨪋\�@��7�[i�$8n���aLÓR����=��'R�D�3&�7���;%T>��Tw�z�(��҅����BIl��2"E&�e���k3�_�j��	K��e��9^~/�櫪>�W�E�����OK�<u�l]�w����6����Ɣݱ�RcZ�y������<E��:JU%���U<�< ���nKG�|��B��A�������  ^�p\ri-���}��	F>���M��2^x�/|3Ũ����`K��!�u;�w\�o�I�!���O��cx��ŗ��0�H_�`�c��+�B��??q��'��'RP6�Z���7��|;&3])����-�	Q�o.��@�-^z���"�֘�2�_�%�吻k]oX��L���7�2��T�Y�wMF��t��z�,���Z���o�H�x��7��� ���� rS$Z::p��� Ȗ��ƤnOa�g�V-�G�y@zgC���b��iZ�P��_�����p���O	E��\?��=f�0��M�3�e"�A��)ǋ��U�u�|�4Q9AE��<:a&���q܂l�Cۀv�y[8�0Ǉ��������ʷ�ڻ?ۆ�����W��S��,;���5�$e�l^���dϱ(sT_��.��zvq�>,]�i��9����ѯ�:	� �%L �8����Z8x������7�\2.,b�qz�z�]��3��!%+��"0�r������`�)ɋ��U��aظ���������u[�ڈ�E�*�p���tϲ�7VVE���5��P8d �R/���@=�ʖ���6x1R�Ht�l���Vs��l���(�KrK�GΊ��s�X�m��I�����l4kP�j�'/)�+IA��Ou�e턃�z�8;�9|]ٙ��$��2LW$8�`J֘�M��Dx��-�b�z������}�7^c�2:� �Z�<��Īd]��l���6x��-ώ������j/�i����5��[X�SR&8T��<�%$Q����K�I�5װj��>����J:���c��v*2�sG𤷧n��f�F[p��D~�E-h?�9�$�`��p9M�㩊^�X�� �1�$DM�7�/����u�>/O��u\�P<�ך�n��Vӓ�l�6�u���4��T*P�_6���P���#}� VSR!e���3�S4"Ē��5��" �Lsٔ���M�$�^8H��K(P�����&�����.��d�B�2"&��x�}�@#8/5RJ����1�ϠDC��jR�/6-F�v�Q\=���˫0g@/�l.Z�E#���oI�1�k^CU����E��`���\ '�W0>{����Ě{����$aIc�mG�h��sk� otɩ_.JB��>�I�M�L�l#�q�7���E?O�[���9����աQ7֧vq�Oeձ�#GH�+kX��Y�`w(�6hL泝K�3�j�m�oF �S�H�?��� �� q�~�x �S^��'��3�%���)��4`�$q9"n���:�0��.r��o#�b�|1�_h�/�]�~���`F��;a�	垌%��ǂ4�Dw�mh���֍io�I응Y&��zv��`�q�Wdۇ�=@�\~�3d�=)�<m2Hܪd%c�ޢ���8�<�z�7*�����d|��G����F����LlOT�?�Dўg��7�i�}��v�I~�����E��ܚ��z'^m�NO(��9���m̈́O���J�J��F�B����3S�T ��l`*`d{�Rl/^>�!���$^�x@��_�¶��)ֈ�Y������H�6�u��A։|�J]_ ��WP�SY?ܒR�a<�GkI1m.�m~;�U��~[�'��f+��7=ӛl/�	M�be��R�[�NG4T��Ha��E�nY����!ا
��*�f*�а�e�&tI��:��'b�I���s|i��؂7�v���P�v8�����������&��)�dI�!��3î�20m(�c'�c	�<ۥq��k�؈B�(�+:lW�vSm�����\��`Q�Y�գ_(WE����C29�@�%��|���䩌��)Y�+zc�G?�˘�u�hN/l�,�A�	�
��V��|�tr:���1�D4��?q5�
k #����P��aB�8@�P#Es ,��t��^��w��Bn�ͥ�ߝ�b���5θs)�mj�U@В����,2߽YT��pIͅ����|23����!��ge?�8�S�Fb2�'�=�n'��+���;�U�����>U<��UD`�����8�0�/�6|F~
*�n�5˖�6��V^4�������gۥ��r������To�;�%q���pq��8��n�^R|��J��Q��oA�5���2�nKzG�8�Ʀ1�$�m|R�3�u�+��
��i��O�G�:,�g�6wB)�[�ݹc� yY�tZ{�P�����L鑵����#���e�(���)���a!�AD_�n�l�^W�| t�81\
��� (��r4��KhMhn,2tJ������w-F�+�j��Q����ƛJ,�dx�����u��$�i�t9�Q��Ϲ��0�����>�������r��`��{�6t����1�_��'��$f��}���eϘ����ʕ1�r�3��zg�N,����㼒��<b�6s�xK�/4���^�FY]��+PB%h ��4pm�4Jj5���w�k)YԐYWK������Pb)?^Bv��-�4�5LTjQs&#��FK���Ž���&����#�	�!X�+v3<c�(-	o��o"��j�e�/c'#y�e����~�d�]]i��H��𞻐c���A�ӕ����'C4P?w>��� -ym]^��O1�����h�:�N������<G�7�1Q�Y�����mZ\j'NbX$^��}[�s����x��7���(DEcN{����N�l'A�FhC��l�Џ�U21\�4iӮF�!F���^�	�n�����M�5��(g�"#��������$���"Z���ΠCGo�G����J��A	!7��=;W3S�]��LZ�ck����C7��g,d2���<s���5t�B�_��`]}���y��B���NJ�]�<p�tx�|w��4�9��UJd�Y¡�%�{_�څ�ij�2��VA�7�'EW�� �&�ߋ�'8{dl�tї��eT(�s��s���T��2�@3��~�j͕�Ni���_��+O��N���2L1�Y���0Q��7��\���x�mB�A
k�K��'�N��)(:�cWKПh�ݾ��\$"7iכ���po�γ����L��n��W���]!�<��"4�|��|Ì*��ׯZ��yX�qfd)@���,n�%\��UL��XF�f�DSvʫ�&w!��RL��R��0j�&���F�ѓ%R�AR�o�1Z;?j�mJt�㭎�A�Q�i�J�m� 8�Ks8�H�b�:0�?�/��W0���u�ĵ��86�2�O�,�)c�<֥`A݇���<�^F����p��j�:'��X#G:�����u��5���С��W�e�T+��D�ޔ��\f�E�Jb��IJ��̭Z�����I~��=G�E��F�m�CP���"���-W�n�oA}P���?q��.�� �X��J����*����Ef[;s�;����l\�`��K׽�߈�_�m���H۟��*�O��CMB���mF�Y����wK]�KY�Ԇ��"��l�R���d\���\F��s�۽�ԫ\J店n����kq�Gy��G�v�-����_`S!_�ݥ���]NZ�C��h��hF�K)�:�ĈhW�	Dp�
���Uo�X�Z�q�e�C�Z%5m#Q��Z�%D^�k�n��(L^��Aa�������޼�F��6-��Φtfr���>2)�,4~JD��<t�,��k.�jSk�� �,���*��1�8�5�Yo5�;���U�#�zw�,]����}s��j�o@�����|���@|�(r�T��E��5(��Г=�W�?��^�_�I�d������8�#(��B'A��ޗ�n373��n�'��&����­vb\[�fg�U2�_�\M��h:^�m��b|ۖ'�.��_�GE��Z���D�hy��������
��q��>M`�Q�t[��v=��ϣ���:���Raf����C���?S�&��z!i=�'}c	ζ�J����ң(4ӌ�*��Ak���_��H k�!G4���8
����F��$5��ʿ�&c*:��K�Q���������խ��Z�L�32*���Bƻa(�Ў$>TW��\�ѝ��)��}u�ѾQS(�D+�t���*dj�����-��h�ĦI��^���2^]������V(��N�L�KB�3v�.��%��F�j�w�&���߶������É�܉c����#k���:�x�1M0�U2�)�7�o�"������5Y��/�L�ˉ2�2q=F@�vm����[���o�W����l��M���M1j�c��^����I#�SY�c�~9Č�j�0�O<�s�'��ГWC���~�l.!�q �7�=�#�o8䍭�@�%�F�13�2�����@����"��_�`���+yU�!�0с�kl��Ұ����&��	�p���RRė(2�+/s�coh�2��{���R(�c�$f��C�.��(A�.G���jŗ����Ტ�n��2z!�|�{����C�r�,����o���c"��`�I]*E�~֢6#{0���5eeI��-�{Z���5o��Z��kNF<TX�Sy��U�B ��iz�ݦǟ_g)9�%K�y�М�=�����q���	�/�L|vF��(g��e�Fr�Vj��Gw`0�����2 
i�.7qm��l�*�pd��j�{#:���Z���S��Ӫ,m��yiL��0.vOdפ ����-'O����}�ػbv`=�h.^��K��A��r�!��Y�0��R8�n���,�~��y:�z���*�W��{���ՉA�<?��!܀���P�<^%t�FI�hdJ��.�?�*���c���Oo�;�{��/�ȫR�a�5�q\�'��@~=����M��JK�tT������}2}'"DTZ�^�CQD��d��壉/����/�𖆓���{=	1^8�U�H�d3<唿��c6����1�17¸jGQ�	���>�`�k6s�E!�iN�˶�r
�p�-O�|����9�H��6j�3i."�L�y��dS$8�
XǬ��(�C�O���.��mQ\t�fKa��D��υ��X(%��A���e��J�����U�8�'2
�ѻ!������ÆUte�IC|UDA2����C^-�<�(u�b� d�4���W���l�$ڢ;�6�_�^@2H�c�ӥ��<%o�c�TBS���tJĢ���3fgNSۢɨ�\�w��p��kL��^�gJ�;����/1*c��M��wTi�/=�ep�ߗ¾�`8��cm�.`�����N��MfV8�}�6�N��񿸏~e���Dt���hL��Q�����e���
뒕*u��Ţ7��3嚍�)I6��L|lN`��T�����ŭ�xN���%`��x|�T�n�U�����������bT��fvx���u~cZߗ�Uf�G��[�}�.�1i��J�$�*�;ߋ��F��2䠇��� �ܛff�2���K��Y��ۣ��>N`F�K�u���dŨ�2o6cl��W�=��* �7�zS�P��u��}�*���%�2XL��8���2�8m��lcLYަ�J��A� )��>���| JFY��3�(��s �|�4X����»ҋ��i�Kx��c���׃�#�~��=�����i}���S�=�g\���(18������CJ�||��n_k�>e�N�R���S+!}��4I#��ڝ�C�\��<��18��޽VB|�wAى{`��S�Wظ�F"���&_G��#pQ�x�l�t���.X�Ń�A��w�'��)��h�.2q5 �۶���h�`�no~h|�ֲ��V�l��m�1����O��b�%g��wssPu��Vf(�[�Bn���NR�"R�.!E�l�<����u����쁡��G3��0��iSS�7;Q4,��wE8�V�c��l�jK��bH�j��h��,JơZ}��\:��0�O~FI�R���b'�I��Qu*;�"��cs���bB&�޺`�VG�?h��d�PH^V�e�ʘ�-�@�V�#;h���}8�; ��ah�W����).b���(�t�bx��È=}}\ɥ�i�a����
|a����;XrY�I�jHl� ��mg�l)��M�Ty19*��ۚuL���&��I<Oǳs�s%1��ۥ���P�sYW�����4,�3����>�'E��Y9�R|R�[f)i�Y�BľğaU���xΓc	A��>,�N"Z�x��^wH6�;0������ܣ���>L�/3���*:�o�=R�Q�`�0�}R�ٺ�$f���O��@�:j㻋F��R�!��7���	�X<����|�G�/���]��~U�L��
�/�/��?�\Xڱ��V�ۚ�q�#R
��k̻zw��:�L�~֣��z�ג�5�����~���oxp[��ޔ�`�	��f�������W>��vT��<���4 n��f�����"��h
���I���cbb=8���H������Q�^���8����z���vf�M|�� Z��Q��Z=Sw�ҽH��l�����AP��E
�n���Y��^
�3ܻs5
�o�>m�Q�5]������n�`Z���@>�/$dt�m�C�w���a �~ɽ�V��	�0׵M�K4C���K{c��(�而�������MX�gQ6��n~����"���
��[0\$�E�������B}[��j��p<%�h�!�Y�@%����f^���^P�@N���qx��wH}$��0���ۈʗ�S�"��d�r�\�= J94hchs~K�i��߬��Tfk�1~���r�������L�
��n޼��cQ$��/~��x�P�D�m�h	�1��-X��d#��)���К�W��z�2~;b���k���=�g�k ��u���TK�HΏ'��� 2Ī��D&'��!.�q��A�uBļ�!��˧��^�t���E��kX�.�F��7*�#���5��=z^Y91�M�����`_���H4-���0i�H�>{}|$A89�
����[�Ln���3�-�XT9��XJ��$s��f�pls;����R��{I��}5,E*�xk����
��?�*!	�a��#�(��1�
d�G[w_H�3o�([f���Γ���Lz]��?E'4����_�8��J��8(����jR?���O�d`UM>w�O��9��{v�)��%�����&?��Nk�����y�M�&paK�v;��f9�%���ʄkEP�O��o����9��W�ߡ!1��Hkad�X�iڹ?�u@�[5Y����� ���.��=k(��S���r4e�L{g�$������Lf���|Q�?Խ��)!Jb j˝~y��;^c-�zN��҃���u�hyj������Ff<��KHJO�F�����n�q^���'��x���]�^Q:S�� �k����z���cW�����Qm㫥R���6�57�
�(ޕ�'�gRN�}-�nKzq�����W{!r���+ߡa��7!�S�� ����#?�=e{%�=]��`�|����w���Lk�'H�6��c��%���I�IF��w��*�����eG%���ѩh��������_$�W4?���w��B�g�9�rH�S�HBn4�fEU&=r�-	�U�Ua����3WjK��2t����l�X��\����W�ZZm����b��e��Nk�Q~���(o���΢��L�IC^�r�E_��1�#|s�q݁��џF�جN��UǒC�BɀI�;v�3�m&���96�A�܄�^������a�Qӎ�V�����_��U������$�?�i;I�'2̢��U�����Y.=��^hU\w]ն�6L�G6�f�E���W�7� m�m�K�`ԏ/�{6�뱤�4���(���6�[INʥxˠ�IR��P�j"4�:K��.���NhUO�//�Y:�����Q�=99���%Bq���������W��ݼj�ւ�g �S�exۖ�ݩGeVp�;p�� xV}j��?�?��#��� �X����Cy)S���w샑���)-�p��W�j�w�y����9�> �/H0���q�w�3���P�.w\.�(��ۄ�ǣ��3��=�%�{���uG'Dk�����.�(A~C�~���L��e�$(e=����$�H�BO��I��Ԟt@��]y��T����e�i?�(�|똨\&�j���dBU&r�D-W��H@:Az�و1�k��U�}5��Ad�2�s>D��F��.�yXpKL�k��k.l�{H�dÀc�p-�~E���S}�)rC�:9I�~�����
d^�jy����a*���b��M�aF�]geڣ���U�^g�JȐ��C����ٳћ��-S�rǲ�.X�~�ґ\
�*�t��O|ސW����?]��A�!iB�$�ď恗�&�m�9�Ur:�E3���ȥ��D�:�%,��_��f!GP����{R�+�o*R��#rC�9��:�:҃����\�*Sd�����r���!�]x&�'扛�Bf4��i3�|ξ�z[5o�n��#\�$*/<�W�cl�#���>!6�n:��^Abn�S�pK����5.'�L� t����Z�ʖ]�ʀ��|A���8�)�WȂ����{ݱs,� R˶o����7Kb�Y�d�?��o4�� ?d{�[�f�O1ˣ�E8� �,+T�!�1� �����Z�Ө}b�,���K����|h��wpv%�d��Pv����*��M�P>��U\þ�t����::u�Q�{���Ix荤�P}��O�kH���-�%)���u��?�d�������������-d��X��* 74Z��͓Ju�W��!%?����8������NcmBt��� /�!�\3��kw�,�70lo��'ۺ&ρy�>�*�A*ߋWG����x���VK�{u�����Zi�6�ek�UQ�Cz<lA=�-���MO]�fà��H�ʽ~��ab4��v�G�ϯ�eM�9�S�v��P,�=N+�F
{�����ftX̿f
�a����9ѡ [H�h�2`O�d��yJ�� �Н��MH�������y����I�;h���O\>Р�-�ly��eM-���xvY��@�C�l��d�A���N���8z�a�$�o��?�>b�j�а�雎Zd�; �H�˶�W\ǜ���hT:���g�{��q�D@�3��.��"Yv�u����CKL�p��krP��	��Ox�ꕖ�|��`^�t��|�n�գ��dv=Md�5�~)ذ��B�9�g���v�1q�滐��Ț����:~$l�Z;e�FSTX3E�n�y�/fʹ��TTd-��PV��m�eo,��[��-<�H��y�t���j?*W�Z�c�&���-��i���6ܸ^�oz��K�ܫh��M���V�/k24�L[��`���W�\�]NŻnz��E�T4H����М���zD�+7QF��Ũs����g�]j�}�z�� �Dh���;��C�.i���Ke<�d	����6r=�v��D��R�� ���_�m)E���㳶�O�(����w� ��yסnǽ�Fd�h�:�&h'�S�����\]<���g�Gl���¼C��9\ v7j�a�~\��s��`<M`XL�A�پK=�( Z��8`��	�䯁���,AFd�|C �[�'���|�뺶Hhw(V��9I���ˇ��N����ϩ��GH�N�,�Uɑ���KT##N"��Q�K�.$3�Ϛ�^�$Zұ������R�UH'�ڄy����|̩X����aA��g|p�f�d4D�6�1w6�
�ޝ����ъ���
�����O���x�%��A�a��*?�dSR,b�p�$��m��\��(���?t���X*4���ǂa�݄o<$D�Z���Aѵ� �(E.Jj�L�S�?¼��Ck3:�glC�Uv�	s�sf{f�xK걞��9�b�Ӽ2SC��A\�n�H�"��?²Y������!K{�$��2v ���^^�"����R4Ϥ47����5$?��/�Lro�x�]N(��&A��/5��J6M���ֹHv�K��n룉8�T�r\��<vf�B z�-��oOI��;T<�M���f)�7j�,Z-�*g�G^t%F ��Ȣ��N���b��թϹm��Ѩ�K�c�.��""����AXrytJە��/�lu�&�Pᐤ�傾O�5%���#���z����	��S�)���3����x^�ȗ�]e���1��͗��iN.E�[��b�bW	�3,
N�}/Y�y'�+IQp0e��-A'cܿ�r4!�|����R�
t��}��/�/��&
��"�>��+3d h�֓|�G:=	y �ʑ[8�{��I!O2�x4���r�#���|���LVʼ��_��Lq7oi��v0��F��t ;v�>��z>|vw8���/�}����Q]�cWs;g�=��
�a�ɐ��?e��Q{=�֊ůjQ���iLB��~U��1��&��q���DMeb��o�$�Z��0N��*�>p~@���)D��q��7�8\�塞����9�:�@�+m�Y�ȅV*wu*᣿����d����aUdQI�����ۯ�>����X_�}ˋ����j��=��( ���wҴ���;պ�W8���Rw`0�+H�02Hɋ��J&����E�#z�I�d�e=u,ם�� �,_�'�
�-H v�m�Q�/�
O�s$������X@�@��Y��=�1�KĀ�
T�Y�?��ry����_',���l;���>����<�6My��|�;%e�֑ 	zM�|n�mxݔ8x/�mɀH��۰�*�;غW+��..�ٮ$���]״�2i�]�zı��
���'��v�(�8��$A��wº�{,�~��r b7����Ћa�1d��#l�j�S�S�*���6:�=}(�i:w�8����4*�?�I�D +����DOaQmU\|�hfhl��qͭj��Md�������*wݶa[)�|��DWz�Hj?�ͻ�P�x���{>@�Z9��G�B����|�	�h31)��}�U q3��u���������qrD&~Rխ�`*�l����������������uV�i*�H�� 6�g�s}�i���"L���w�	q���fm�[a\�;���R�|��3�j�X�vt����6A/���-I��������V���{�F\LAG���ɅIi0<i����6!iT��?@�lU2T�Թ��P{B��u+R�b��}:�24
�>��)�vr��ܗP�-�	 5��	��p<�/�����B�3�e����s�$��X���'W��9�2�� �`�<5(�`��ۜ��ډ�|���k<�1�w"G�t�7��l�����!�_}�5Z����c7�K��Ĭ���%)�������rSMӤ/T��w���P��^l���j�O"��}!m�ɔ����U���s�j'AE��iGQ-�j�f�zbb���9���4����i�k<6k�F��k�o�]��߱�+}=�==TǮt"�����y�d2�~qr��>�yf`�!�K�<V${�p�[z���^ ���4�lТ ���� �4(�Zw�,�Ҍ�g1��,j��G�s5��"����]1Y����bǫ�F�/��T��`��O�$\;��sf�|�&!�_����L��:d=�G��/��X�<�L�C������t��ޥ쇟�g��H��%�1d������ݕ�a�Ժ��)ez��#������oK���lڈ��k�����H1����m&~V���j+%�;��P�** �Ϋ]CSJ���P� VrV���r�P��c=U���������
|/B~{��GY�t���0qT�����&��r���"E����4k��ȁ�����e_���#;c����<�&�p�$1�h�� �ZvqJ�sYdo� ��}��ym)T������:ȷ�
�pO�JH�9�e����[�����Ov9S;'�?���"��cb�(��,�DS?#��}[��D1zw�Ϭ�{I�q��b���Ԙ��
Q�^�x�Z=�����Dg�]:�vkHy՞�Ew��c�G�k���+(��{�N�+`�>��A���z�-	ƶ\��M2��s��m�a1��u�~T�[Є�|��yJ\��s�����Z�y�z�L��R�񾭸��O��XS&]?^�0�<�̇HR�MW7i�qA�[��!�L���W�J��ˈa���q1��![L�i��,BDuk��>bt �5�Thϛ�3�x8Ƶ��YX�[�"�rN�2�1Qz�P��HÅ�5m)�^��R����qb0wz�Ͽ�x�뱤!,�8�W&4W������_5��@6�8�o7R<��>O��TCl�([(��g4x��U�\0V�{ Xv��+�q�`�����G����M��K!c��zO�>4��A��y���x� �1�&'p�g�x��M0�� 8���B�`�b
L�4e=+v[���ͧ#פ��e{w���+�F4��qҥ�ӭ����Z�Hc⼈��l:���zD=�X���B=Ҏ�����X��J�dp��sr�����ಜ��g����C�Z��� �z4D��i��àԠ���,B���bk�V�&[��+{A�)ϒd-|���~>s���r֧m��l��m����޶Ux��\}��ˊ��d��Q!��
� �Z�c� �f;�7�r�Qh�{�s<p�|~�KB���wJ��i@q�R��'1Y�
��9����;g�R����s ���7{�S�����KhD�5��JP~�a�{�a$Pg����;z1�>I���Xa��H������3OĔ�����gzV|լ������$:��}>�L�U�Vq�Aen_�۟�ч�٩�i]H��\_q�+'����.�K_�nZ����ө",��_���+/�۹`�N}q8b1 �Re�v^�\y�%�m	�)w@���<�,�/����9C~�->��-�:�K+�%����;`�by5�ɬ�K��A!h%o��%}9����'5�߁>a�Rp���<=k�Mz�1ѷB�	�b�(���d>��yG���B��K�')� �R�RXo
b�m��h(�H���F&2�n���I'k��j2؍�Ќ�����sX��NbU�O�%���-c�_i$���I��E̊#$i����/�W�8|쾶ǻ;����9�Am��1�w3`�_$�^c��g$Lw�s��f2�Ώ�W�6��3μ�ox:!���0NW	0#�{���nd��׾��YL���z�r��1��G�Na�#���+Fg��������ƁF�/�o��M��KP���p"���D�ą93�Ue<�NZ>���P3޵�翬�?�xɋ���х,8}m	����d�jUtTr[�<�}X��q���*�[L�wW��h�2[r�N ��FMm_�����E�t'��"(R��qR�1��vL������V4�K:l,j�/׳���s���0��XH�|�����:(�+m����*�`L0��y��a�0r��cT�k�b�r�����D��]�(�tD��Qb9blD���Ӹ��T�Q<ฉ��w�駷B��Zn~��q�gh�6GEr��v{Y<���FDzd��`S���zwu7 a����x$�Q=k�O�{C�ϩ��F-d>�� �OU����u�QJt�Yc�P�LL���!F��L�i��S�}���4j���m̒��P���e��OM�
�h�3s���	����^��Yg/{[C8~��D��YKȷ�X���>#T�����grfA�LR�o
��g�P>�(��n`F�8��&K]���{Xĺ�a�֧V��A���Y��'^���8��z�R2���$Tbn;�f,����:�=�6��Ē���GKTڂ�����T�o�\�_��X|���� >�e'F'��q��5b�p'f���[.x�a�]d#DO�-���-��� �a��4��E �ѻ�ᾉ�g�M`�6h ���~ +�i{�p��"�b��=#^��W,WJ��Y���_+�΍�#%�saQ������U�Чz�\���
v�����[Cj ��8d�-hR�=��e.ݳ�&_��Qf����33���#M�VxzJ�)|J�/mS��]�nE�r��Ѐ)��Ka���3��<U7���o�c<�YE--Mee�0�W5>s��9�4��&�7��-� m� �5����}�!�%��5X�e��du��A��ʢ���ئ���TJ
������%��g�޻ٗ��њI{����K�����*O5���Zuzh�������je��q���c��4�j��D������=�jV8%�jb��Q��,r�!�չ�^�۴YW��b�TL�{��?�=���"�7��2&*4�	�����ִ�`�N�$D?I��B�e�wHb괷n!�%���^z@S��>�?���L�"Rq o��|f�#}�V� .�I������T����\|�"��_�0� �����C�����)��"V�h��8�Fմ�Kn����u=�yO۹*R��`$9�\X�z��&d�Ωm��1�]��6�$�9�p����߁|u�����f+X��K�(	V�qL���h�	���z�}�	yŠ�3�m���U) x��*vٝ��4Q=���JR��<��4���z����d�~��w�۹qP0�s��C7f:Iu`B����K��g~�����i`�d��(-��L���(��C6����'�SK� ����'@�s"_�Vi">3~�����pW��q�wK}y5��������cK���O�T,<�]N5X���G���k��Y�P\ɾ	6�� �9�)=���Z�t�zc��r2�@��X�.����8G�NX���/К*](�S�Ʊ�>�� 8ѐ"��Q@��Ev��9(�>��`!�$Ԙ�/�����M��N�`�/hq����R�R��8S��M	)
N�X3|�h?��6�JE̝kI}H�;�:�����_S�CfКe�W-�zk�}9� ��;sD)k�	X��٫7@
�l�J��s�M�l��u�dD�{0_X�#���pzc^/�WR�(�<S?�� 2d�J��8 ��J u���t�n3����|��>vҐ��-�(_�=1���ҊwGo�d!�/�ڥ��s�������nrؔ�����y!	�S� �oR�ͽ���kqҲӂ�T�+d�o��<�_�2�7KY�xB|�L�L��!�'؟r�ntW,vvp� ��+���y����� ����%��!���G��&H�5��i;�j�/�y%T5�P�I�b$[@�_���&�W�����bז�(��t]��s]�� 1?�s�^EG Sc~UX�K�!fh�K��<�v���p�=fwP��$/\� /���F��"t����&qH/A,7U6ϲg��1����.�Mʆ����֌��];�w��f҉�[Ӳ�&��������� !�_�l��3֧-��m�*|O�!����W���}"y�0lʫ����]�ԭ�G�ϯݡ��E,�Ǝ
}�;ٴ W\�f:lflZ��[q�v��D*��2�Wkg�H~�B�<d������ 5A�4A�r!�Q}�_���_����uC�������,f�- �㷻�|mX��ձ�a����3Ue=�r�E���2s8M�L�$e���i�rc�\v���A�J�(�'ٙ7����B6r��#��6f$;K�HZ�ZxK�����v-�	�Y-q��RL�G�����ͤ�t)��7]��cS�H��<���DXB�n�|�F�o.�p��h��p�ҬuH�뮞��7�sI�������R�FsK����"�O�R\,���-�/Z���.�P�?0��G��t����J�oy	괻2��x��*�:�l%4��?()����*�*�
�h[꼇�~�5��g�t�9NT�Ϙ��;:I�$H�3r����?�uM����l\=��>�:_�f��A��I\�VJ��I��%�I�s��`���;������o`�iƴ�ċ9�(��"�� r�W��s�k
f_u���O�R�zH�X�g�R�VVc��$�f��n���S�®�:�qn^��Ȫ�%ם{�3�(�2��QW��2��w50��D�Z<��J���T>n�'"�K���6��JvGGC��Zܘ���%m�ec�w`s��ܺ[yC?�>�����.R2(��5ĺC��+M����s����|�ZA�`3q<lb{�[��B�ε�)��9X8��ӂU�0�^
�Ԅ��w�a�*�h���B�+�{{�c����i^.��;'Q^3�,7�[^GQ���rwLH�DLmѰ��P���P�"C�u�/6��Z����?�/�uVЍ9��ď�EQz39�|t�=�[�SmmdI�`�h57@��Bՙ"#�ˬ��?fB.�ݪ�M���U�%�5����iT Y��
�(������b�滭�6�]�*��?T����s��-�zZ���UXx����+7rM��T"xW	��K�_�В�1�����V���Vy�Cv��{BQ�Ԙz�>���֖UN�Z�yvl�E8��=�-�����H��ͮ�*�*��A�s�Zç�0�k���8�P�h�!cSje�����73ս|"�M3,Y�߉�T�ﺽ�5㷈p}� ا��?�w�B�dY�'�\v�ws�Et9M���ݳ���y�C���F��
�{�]*ٷ��r���=�qt����_������nލi|��P�\���Aj�V�D��1��`f��H�F��ݒ���5,��b��l)зB�� xԩѠՅiJV�r�r�k�L4c2�L	�J\i/���U�ҕ���J>��6���1�������e%�9�^ѝ�-D�g��Ԑ0<*Êe#�%S�aT�R������q�%͋Pi�-�o�a�/1�P���6��_#�u~\�@1���eJ2@�{��7 �Lw!��9�lhL1�JUp�b:�4J4Qh��7Dt�K��%�>�s�9��t�-UDl��(8��Y��ZR��Mb�;�����x�|\�]w�ɠjXYo<a���﹀QR\s��s�3u}:���,�I%O��~�����!�|0�4����tZ%���;N�:��a�'M�\�sd��Zv׸d�"�{��M'<���I�+W��h2��}���{0N���ɀB<�s���C��V�W<����\���u�w�҃��\A�|��'���~��R�x���Y�A�	�
�܅S����1�lI&�g��H!Ӫ�f�#@s�]^YA\2.U��p�D��ʘ���;��oM����QtEuLL�t����lL�\y�E�hZ��]KHPě�A譫�P����K�2�W!�b��qҳ�/B�Q`��D�YۮX3�S�#��>���tWAq�Őo4���E�@���2�����1ځS#|�7�R���/��ي����K��ʦ: 3ztQ��*<�س�����1�����O�\Т�O�u�_�F��ms�����hu��A����Ml��گ�ņ
|�rNlS� tݞ�5q�0��5 'HV5���!�������K�ΑX���w��- ��DW� =��o'x�!|e0���ڷ�槵���Z�\p輯�·v -�U�e�}��{�����ޛ?�'jJm�
��U�K�<rl=�[_��\��H���4�8锕՗�
F:\8 ����p�OSZ�UzC��Ce\S�'�ݗC �����Uˎ�-���>U���T���m�k)$M_����p�[���H�dJN�=j�,F{qӭ���� �/P��Z��*I�e��VH����h��E0���� �$���s�b����UcZ;�ZJ�����(F���P����ZAS���-Q��� ��"	�� �I}�" �4w�Iv��l�-i��Y�ټ��P^�,�b/�\�W��|Z/G:Щb���0�Օd���6�QV�V��t��McN�N�uї�R-�ᾥ�{1W�5�pk�Á���Aq����>�{Z�1KF��T{��;��蓾�IA2p푅-�D	��z ~&�ilf��<wN��\��ƨ�Z��@ly��Vp�Tpp.�ud�͸�rϺ)���������u�b�]���8G��p��4��mMAWNt�#�4�!�2�Bf@	 ��u�����9��$'����o���Ӧ����l����8}�R��=�p�ZjAL5�Dp�8]s��ku:���:/��~���&��^�?�e�ٵ���ݤ�.R�5�Y��$�0�;���Osgm����dq���J�̋�5�b��&dz��"��J�ɨm�i�3��[�ʑ��;�ʃf�1�L�ǉ�h�I ��P#jnP�V��f�/�D�$ׯ.���o�������QY��V�}�T�q��Y��x<7���
Һ��?�Z������+ڱ���M4�yJ/J=U�`�3��Hg F��g�8t*^�ߕy��?�կh=}�p�P�e#s��7�:&m�|q�hp �/Z^5�-vo{#�@� ��P�aqn��g�ަ�.ޯC}R��Q/��ҰV��/��9 Nwm$'�|<�Er�^*�$��M�S��*�߿ Nņu��`W���oV;����겶9���O�o�H�	1#k;Yz@]!�A��n����f1:l��n�ˆdX�/8��V�+��NB_�s�·&�4�(Z�t��ԥ���i ���^ �
��M/Dv{� �z�˴�Dr��y��{m���9cd�ʥ�����bP�+c�ÔR�x4>��6I��-��(�-0(vA� B�_��v�v �?Ku�|����e��"Eh��Ewh��;����)�����ͩo[�*�R}���Q*��n�F��\�oW��=�A^\�}�׉���IN�jNK��,;�nq�F��E�=�gkj�K�#�y�m�Ӽ�(ς�gu��l��U�#��o@l)*��$�ɿ:$����)��=��6�[��qUS]�� L5s��Z�&p��P�&<+10ĵ�B��ȅ7;�SS�����Z��<�(+��zn_k�Pc���>Cs-*�~�a
Z@��1x�!�m�;d\gTU�̻��V��B�{����\��^�[}�)���o��U�8�(?@��oN���bDs"�u��	��%��W���`N>�]����,���0q�YDUs3���}��7%��6I��iĬl��2FP�[~���y�5�q�04������hU���(��/^�8<Ic�W6Y�ȥ�������n?����J;�-6D0�~ꬒ��am61��dscQ���Cn{��6T#y>!�k�>�F�\��A�Xe�ۙ��^�h~�]�ν����Ù����&ľYjٷ�f �ju큯/ϻ�HŝhNjw]�nЭ1��ZkAa�7�d
۵!H���A�v���5�h/
����G{OΕ�Ɵ���n�	K����$��,�i�7�o��vR�(�ȟ��>����VS<�{�o��C�x�N��1��"< �{I�F�;�r,�8�6�t�ϓ~\/��{�����0T�"�xa�NiU�ɢ�S܈x?�;	]��$/���[�k}E���u]:�>�T����qJLHŽ"NK��z��R^�� ��3���Քi��h;Į�~.J�B�ͫE��=a�[BU�Ԯ��p��Fz�AI��T/B4U< �h�MQ������e�<� ��ۼi�s U
�K�+`���ř4�x�Ff���c��@!�@^N���.��A]��}���� �Z��-m&�ak3\�GPC�}�(>�-�+x�#��h����e@O�+�+��~��ݿKXpB�n=�y�{r[	t����Hc�������[����g9��4'A�!�QΟJR��'Bm-V����%�y��=}�W��;tws��g,����,.��UH�,"�C|����Pɲ�g�ٍ?E ,�t�_��[��)5sw�RQ�[�W��Q���q^�u݅% ���F�_%gp�n��
�jeǗ	�1����SW@>��`)� 
�Ù�M�7r@�;F��'�xm��7�c�9�i$�_)Z��߯	��w6:�v�j��v��-���	���j�)��R�`5�&�
p��9����1�Ԁp喟�G�5���ضY��L�*�:h#�ٻ�.b�t��9��^g���v�D Z��o�yf�#ɚ�Nh��_:/�4���8*]닧k$�j�Z�W*�g�%9K�a};~�B�`=�ε�]c3�N�}��������(����c��XE}�Z�o
 '��W�k���8�������]�a1�b�����bp�F�������Ă������5��X�>��00j�1���{�[�T�jW������2�D����A-��K��,Íx'�{g�i� i�^��}�V�9��`�$`�VF�+/R!9c�עϟՏ�2����;Z�%���4�#�d��}���y:�-tEOg�����pk�-*�����/3�lףe�������ېN��C#b�o)+�>f�k�~�,��d�;Y�7n a���Ϛ�,#УOe.�Y67<����k�$C΋�K5�;6�?��B�xX�k�i������XXC9t�֏�o�@�v,y6mn��ʻdvu��aou�Ҏ�&��=#4��G�]2�6�����-�Q�Ej�F���n�ݩ�X�Q�݃�h�����i	.��oŒ���=���򮳿	e'w��)g�cΗ���9���*� X���q ��UK���+L]U���PS!��%)�^���֑��o��n�.���f<�mY��'�H��'o�X9�u0(��NU��/���$!��EF�O��o�x��4�z��x������S'����>^��vK��n;�����[Bmn+^F\M��n�]=;��=�F����z\ >S=�
;��>X��(NY������%s3{��]c�����̄+l"�~�	d��O?J*j��%ZhN�*�^!!f���RA��4.iͿr.�E
D\A��]�Ǳ=X.i.w!J	�z���ŋ=��( �����&8����o5� t�ΰ��&���o�5G;Z˒���K��t���	8�W��d��qs&H\B D�c���D/1p�˟���O��+P�����@�QY���GJ����R�s��I��1�#�������Vyy$�qQ��_ߏ�X�tĄ�2�վF�]�*N�+���'7c&��*,r��]��nRXt�k6N�7߾ه{�'�?؜��n��?3��d��! �w����e�V�K�-X����v�)��lq�H[p��Sb�Yk�?�
,+S�[���w�ξ�/W�e	\d�
�CL4�E�9�4�	� 䫳Gl��>{UT�4�Mꭄ�q&���ؽzCY8�7h����?�����zh�)Y��'D�q�0�sL�a�i��+e?�t+d�7��σ�|L{5g�y/O�@��_$ ��{k�yCO��p�w�Hñ��m����U����Ky�����Tn⼂������49z�s���HuKY~^�Ǆ��~�1P��D���u��NJk^²�\х.�=����f��ݐ�>�������H��s ��%:�VJ��A�"y�>����rZM�2,P�	u �T�eG�}+(�����bq�99ٝ�
���}� �]S�YK�V;ay��H��@�l{�X�Me�>��z���2����A<�H�\u�'2++Wf��Y��bm�^�ŝvz��(�j�ۻJ��o�j�����m��4�3q�{v�8f�J9GV� yn�8��5j����\�\E���h˫�x��2m)$
�k��[h	R��g�f�����eU�YM$��d��&��?Q�i�J���Tִ�<eK�w��mV�k��]�IY�g��}�L�&�PX���մc+'�p��ȶ���ּo`��%��7��}/����㭘wЪ 
� �#�/�2��0�AR�v�]��M�jy��h���{|	*.���;�R��Û�灈|'�@:_|��(vh�n�5['����3bY-�-����\��c���E��w�^�Z<H�E��{Y{s6%�\��e��8>���ё4Չˏ��.�a�	�4s�?�^XN���k�Z'�^lF�����&D�}�,�Q��<rkb�ד�Dq3|=�3�b��ǆeB㒾���KD�:PwpP]�h� c��M])ߒV�t������=�L�h��%h&����)���'�s�&�W)q�\���4�j9��ẅ���LE���X�J.&�1��gs�}��C��n�����su�fmo"}ѴV�����45���|������6X��i@V,�K�k����m�3]��e��Ǹ~�4#�A#D�B*�2t]|�J��D�&e�71��#�T�n�lB�v�p>�&�* �Y�t����A���=vκ�K�9�jǑm�=�|_�~�'��+B2ҙTg!4���Ȟ�2�b�T���G%��1N�4ճ�<�	,����gۯp7Eᛚ�xˤ��^�5H�yI f���"KwՊ����ٴ����݅|&���<4���+坭�eG5ߞHoGNN=�H��#�h��Y�C3J10�y��\�]�l,16e��H&�iԵZ?�gv����ezmz����=��DњUie�t��X�R��"�ܷ�G�Y���	d���R)P��ǥ��@�n6ao?BG�xt��'��G�
h�Ԓ���7!��^S$?X�����d[¹�&�����uD8W����<�T^��;d�2���p"����%T�u�9��:nA�dȫ�믬��T����`��(����E��Fs�?Зca8��t�$2��A����k��)�O�M��``ke'b]=S�^y��D�M�{d�XL@��G;����?�b= ���ȃuJ���$"������-��n1寒Gg�x��q�gUڷ�c�]�<�{荛�3�PQU�z��]QKZ+��}|�^��]�ړ��0��rM�X��J����-7_�����A���@7L��n��w-y��T:���U1�r��yͣ�;�/
*˷q�v/�Cˌ���#s��c������-nz7�������E ��ǌeT� P8�,���}�!��%��]z�y-�������b�۔HYi��?������\�����Hw��w{�/�)�'&��q���Z���"�N0�Ю��䃱
a� x_

��D�_b0��N@3��V�;s룅=��	x̄2K�u��<���9���A�h}+µ��_�����Ԙ�D$� ,�Y���T�
	\&%ƪ�)y���P�Q����*���=N�#d1c�0�1Ծ�0$�Đ�R��`ܯ�OP�M<1,�y� ��~�ء�z"M^{T������t�9�`�P�|�Y�<���/�D]����k9������4��v��rZ�	⣥E����/�Dk&��&�Ħ�.���y�Tgk����:��ZA5��>c}��9՝Iϸ��P��(#wKkN�b�g��Su���)&̄�T�ؚd:��A�ڔR��h�g˵;�S�a�ηm
�L�@�O�` �l�F~���e�9��.?k����^���+�Q�)& �vX�aG�_�1�#<T?^N�?#��2x�e��L�9�:f�:6'}4ə^;�)������=R(�s���x�@�s�4Q�
JFs�=�5A��7u�J%f��_�m�����1�i&9x���x�w���rp��Н�j
�V�5q������i�9D�Zj�D���H���cR��C^@��*! ʠNG�t��4��E�SP���3||�A����k��P�,Yr1���쥴ڵ]�Gh-}R����\�dAteX	;��\�s0x���Q�U������}���cƝ��<T1��f�VC`=�,|����,��6H�2�qS�X"X.��]=	�a4���*(�r�BZ�K�6v\MF��� �f�16����d}��3!���%�V�����Y�`c+��<r����$���ɕG�R�a)</�- *��J�#�U�e�Z;���:y'�+���(��+&�<�NrXe*�my'F%4<���i��![�yCȪ��2sA���%�!���&��;�fC�+D6��NJ|]�2[�sf�L)Q�q�1���k��
Z�?���͛����V@�W��ђ������֔��c/���`dk����~Zu)?m"lzp 3k�@7ғ�Goz`�����!_���*D��q�y\��2T+�荐QHV�k�wh2s$��`n����a�%��>Kfفl�!�I����NA`'(� ;`�g9"3��C{-�k0����R�d�R�@T��YD
1Ng0u��;y%�ِS�ML�֢�w*-Ռ��FW�^�
%,2Qi/Bp��d��=v�K��yNG��?��(�JNf��[(����2�6r�S�&,
d|�绿����z��97����.lȘ���2��[�AlRsw��䎂��H9��}9��Z�O���9��%Pr�m(�m��d�U;m4g+"c%ߎQb �*�dYjW\�\��elݖ�N^��#�L6����{���>�\�5
[�s��Sׯ��?i�����s��3{���N�i:[FRJ��E��������CҼR����1��&��N�f�B�ј�iK����;x]�ۦ�im��*�|��ȩ%�Ҙ{��N�EG'����<Q�z0�&!tsJl!�i�#mo�6d�}��/UdW�鿤0#�+8ٶ���x,�Z����
�&U���8`q��3s�8n����[㉇(y��ʆ�fy�m&3���ujcŽ�����I��p�;	׭U���:�!J���%t��9��F���},��8�RK�;�i��%C�57C�W���1����3��XW�O4z���-Ǔ���~�(�6Wo<T/t\�t��?/�\���C���݁�������3%;��M�����9N;�E�g��eV�*� m]V!�~��)���J��EJ�Cl+x�<�#�!�a��S�ΉKZ�Oy���c�&8M&�M�қ��ʒ-",�(�a�l�R	9l���⪦n)��(��///����`���9N�Tw9,k�<? P�\v����)�u��x��Q�!��m=��3�A�T�3*� 	��]&74���G��%SO+rP|%��B,�*�t`�����S��Axw�̯fg$��j�N�_٫��3����?��'�i�p+�O����s{¡
�@�������`c�Y�Ş���ѾN��w�%Q�rW������d�~�4���þ3���M����5N��Dnt�f�8�a�~�ys S���Z���#V��/{"��Wf���A^����:�4dM��5G+֦�\�#;�Ks�Mj��!�l�)�~1[���*0ǖ����	Z H[��L�m9,tɬ����C_�(�iB���H\|��W��}��9�Ʊ�}VP{O�ޞ��j���O��\����fc�zBnP=��w<o�c$�1z1pl�H���|�!4���H�����s?9v*��k�(I��ڐT9b�Ϙ�LD�6{�_�O�f�]���{y��#�4�dB�:�rg�S���'�W�f>'��Oŏ�L������} _���]GwGm��BR^��h45��Q�b].<���+�4�l����`��x?bP��R*����'�z	p��Ŧ�%o�_���J�V��h����Y�������9�1�>L��?f8M�t�f�������s�XF��l6F�5cq#A�eK��\Ο�S/ ���W�
1NO��i˩�,e�Z/pE�勡h�,��s��6�H�R��Z���dR�0�q��_��w�ѥ~t>�?��u��0��;��rg��X�&��+�@��0��]�O0�	�m�%/�ݿ���n��V���?jBG͝��.;��7�˄��|D�O6�!/[�+\��~:��u�7x�����w+�}��^�'-���Ǖ:(��/��d9���6��P[_�.��P�@�4-��la��)�~j�g�89|�D�a���"�����6�+�B�X�R��*�f�Q4��f���p IQ �P�R��u{���Y]�e�Q��<��+�&l����lP]����ۿ>B	��A�C�aS�d���o�+�^u����mĴ�����.�<�RN��ͬ6}�"@�T�D
�rF�U�����%*]��`w���牣�z�T�#��9M�r.PQB���B�c��x��R��p��M�Dk��������3�_pl�|,�ǎ�$IDʂ�"��=`�.0���s��n�R���-��O����0M�\w`4i�8�A��H%�d��/��g7c�!�5�?u�P�e��B�S���PN;g�- ��:��$����]�rG5*`�{9���S��>'�	�t�bs@R>$���@է�������O����äX��7�*U� BX���'����#�o2�~@���n�Sa�3��&�\-�2 �\�ֻ��3���T���㎸�E�UJ�scC婱h�f�T�?�%4�=�.�'��t�D���_'09_�i��9[AT�x�)�u����xP�q����+��
G��Ғ���'z�����p4��,�x�F����6Bi�{[����K+��v��3X*#B֎�i����m�:)�B�����*%%�ҩ�eSY<�5]�B�r N�q�SWR�_����dL�_���Q@Z�p(���y����"�^��O4���٫po�u��'���͙��K��3�|hU��bovׯ1���Y�$=�Dt��Q���j�u�%-Ό0(]f�9Ve�c���#�����F&�F]��󢿉����JL�h֚(�������3�C�ee�j�<&�G�F�<�m�j���g�h�Xp�8b>����΁/��o���O�VO���KH�}�@���Sҙ�����$�ļ�J���P����|N��eތ�����i_9 �ݻ����<)���,��>$I��
<?K�y�K�Ju�1�������՚���V���p�O�&�_�<R��O�Y��i�ݗ�?\D�q|g�w��J��&�����X����3�ɸ�5��F��*s�O��bmwU�:�f@26G�m{#*$W4��~��|`�Y$�Ԡ]n+�qo�k_Ar�Y�#�ޞ[��[Ŷm�p9'�Ow�at �����}��G���"J����K��֋�y��Q��y�]բA� p>8亮ɽc�c����2��|��k���_6u�`�5y"�V��	�nJ%!�#� R��U���Bf��m�^��L�
���/4�zkI������X���i+�o�)��v�L����ĲaDnC��Ӊ��� �7G�W|�[�]������ӏ_�E*�_I�[����E,Ng���/��|�O5���-�����w�������q�ϩI�%D����3�Of��a���R��\�ʼ�D����k��>�Ʈvk�RK�Y[�[��j��)����j�6�e�5=��5���*j2�t&v6�[��2����P��j��R��(�3���|�L� ��9Ӽ�!��J����@����E@]�N�p���L�����r��ZMK��½�*��Onu�R.ߴZ���܄u�f�׃~<"�W�=u.���� ����.����2�YǃシMu�]�v�{Ja����u"�"3��F�T4�P	��Î���,����\�{O@Ys�i�G�e�c��~p��>뛯����
r�ggT�K-]���}[�%zO��V���0�o��n��.��nr�2ð����/��Z�Rh�ZǱ�Ϩ����EXl3 U�Y����p�o_i�rE^�:��sͻ���Z�ž�� EQ[c��A���Ґ6w���X	P��+�ɤ:��ً��=]��%@�������7{y��ˮ�;(��)!J�|�0���u��ׅ� �mF��Ͼ�k�&L���%���磐�FM�-�Uk(U� z��P�r�˿� ��^��w/�!b�����Y���U�����Vy[�a�Zy�e.3�G�m [��� TmR��/�����h�B�U�j��Q�4�a|׆"%��)�E����8o$7���Oe����WE��8trP�H{�E$%�'k���W�%�z��63�پ `\�����s0�NqҀG���߳�2M����*&�]E�����8��ZC?f�m��{� >DT��	�E/FQ�RO̯�����ȂWA�41��sE�&$-xm%'#m�q)�tc�����,�õ"��MNtu�Z
��ӗ �C�{Q%&)�#��S�No�?ѭ^��I��v0�:�T���_�돂ieI>������jH�q��r��2~���U(�)�[��=gh�kJ8��n�ֆ�"fV_'G��6|ܒo�1K��Yoa���	-#�,��7I�>�Vmk���{��,O÷�I�Vt@1�(��ʣT$�8�o���doJ�iп��qi|�:�%�1~�a\Q�ۏ�X9�H�����F�$x�R��� �տ5V@��}��1;���W_���v�=]�B+\*���B���_Z�@���qtB�Sy��lQ/p��8x����;g����j7k ���wBoRB��cJ����� *)�L�-P��?"�y�@Gݴ�&/\��7X��A ���v{��oI� ߰>�}�œ���a�Ek����^V(l=څt��	�cn'��@J+�����LO���s����&o��*q������ZUP��֜B���ٜ.,�@��W�N3��[�J��� �0[��,̴B���CE�Z��,�N z����
�����d݉��»>�֠�a����`g�iJ�	���*�����2�"}�)n�(sm�jL�Ԛ$42BF.{<��E*`z�����]���t8X	?�<�$� �S�R��_U�����`�k���y��f��@�qZ��8�.��P���܋urP>�1H �&�����`��"�b<��R3���D%�up=o�Z��O��(�M*m���b�
n��[|�M,�*$\d��v�i'��&�v���X����r���� ��B�G@���hs�O#��Ądl9cc	Y��å���ю��5�
���T8+��<��2ʵ�Vo��4g�˴G^19������C���]����"(��'w�I�#�.f�����b?�)���[կ�4MR��T�,���T���?�-�z�ϵ�iW�Et�^�`��1��J!���
�\6\�N좷x�w�ع.w+�)�5R}d�z�A;�U`��x�~�Aр�X�B�R��T^ɛŸ���k�gyZA���~�u%�q|��lpˮH@����r���%vV�� ���W�\�I�z%].�*�:���z?��|W��LAy��)��.īH�x��U��vH��:�p_�JgP$~�]H�Y����enSR��n��<p���PA�B�x�t��*W����� ĵ5�TM������%�W�X�Xa	�@�&\HVH�*���c(�;])���t�]@�/'c��7���va���R+� �5�nj���%/��j�3?u��I�S&!O����J���j���]�D(�����B!F�Bz��zO����6��:��ɋ�����w���g�M7�~�3�`f|'������/�.{�jYsx�:8ӋEO|� 3�U(�)}gE3��Y�Z���bp�V��?�o7�r�p�#��/�\)���L\�!W,�P��cZ�u����C�h�*�V�3�Z-��G�|�F�~M�}V{G��Io	d͍r�@�,��CR�+�6�µaB(�p�s�Rk�j��<�Eր��Er���6��yQ�Yq��3�N�O�Y����Q+$ �:�$��ޑ�%C�m�U}�*���AE������T� �dt�.���sL�2�<*��?:3em��ƍҽ4��Thm!c���\�t��@ѵ/�#5��\!�;��w7���&٭a�9�~�j3��!��N��v�����	B��L�h��3��C9 ;�PE���sO +�~C�Nx��\�1�?HqA|��<+ji����N��?�Q/��q�W2s�Wg���1�J�A��5E<�d��i���@U��1^�#r�Q�|�$�Ȥ�.�qTo��96��ã���'Lk�\e)�|(-��>#�5 P~/R�ms IkLNU�7Ę��|�R]�¼wG�Ӥ��a�)F58q�V�t�kMb��@dI��oLp	��Y�(x-���[��F����w9"�
%�J�	��{`Yʬ�#ދ�d��.��g��{�<�-}9���9t)�-�vf�}$�����pvTv{Q�)�C�9O�.ݣ�S	<sPŪKZ��9�P���
�,��� AJe�^�����@��n7ٯ��m�"^��RƘ����[�%�ěiam�[�b�W;���>Xէ���o{���=��1�E��0�wA�r��.�s��X����������Sű6��oq���c�Ӂ���Hsl�&A�߰�����y@�I���b��3���2ȳ�Fck�(wMߌ  O^�f������㍢��]�W_��ɾ_���Ww��B���x=�=� r�-�e�oJ�u"������SʤB��a���$���_#���Ҁw���NQÒNr�o+B�O�ʖ�y�:��HF�>���Qܯ�0[�.4>��7����>ސ	!��< du��eڸ,�,�s��a�c}-��"�`�1y�Q����"2���x�id��c�c���8�.��z��>���y�:衅�~@t>�,�PV�a��A��t7<��%���P����C�LJ���+�f�t��I����V����6�E���33���)n�w��{~[�f�� 4T�g��2i��[�n�(�@�����cTAI�l�[�W�L4��%9އ��<҈^���"My[%^��α!-�c��&{���n��ښ*�?��d�T�S_D�10֫�����]o#�n�������K|W�_sY��'^�ޜĢshƈ:�j��nÇ+�#,��œD�8��d I�n�3:JiUtm������J誔=Ί�e�X�����/Z��1w?��9LT�y��ٗ��d�fĘ�zz����v-���P��?��ه��v-�k�S0R�i!Z\�B]ǲ��@?�����^�+�ƥY1���Yf���u����*����?q�3҈Z̦e���-���-��3�)#_�]F��8��;�u��#��E< E��uC�H^Yˇ��n:"�h�bq���l{��`{4�aԴ �('�sAkR�"�mf8��%�׊-��y�u����Ʃ
�~�p@���i��^Ys����a�mgޱFڐ���A�G�HzD:1�~�[�QnJ�^�EZb�F��ӑ�ְ9L���p?�}�_Z1<�ђ6舓$���XZ8�j��9�l+�p^!�~Z]��9s oL��WP�=��M�_Aۂ���Ʌ[=�)fĕ@��nZ2�n}���.1��1oF��y~�Y�uRM�.�U�8�p�n��@��?߿a ���Jp��&�o4��IG��\�{�q�:h%���_ϡzї��F��`�}���|��[5;oQ����c��c�-�o�����d|P�pg N�F|Q�uc׉�#k:b����N�����5#�� �u��ZUl?˹>�����'h���L���J��A)� ��6
����˛^��G�iÙ��R����&��}���N�X#�=}�T@�e���t��l�� V�ݺ�c�n/X��=2�������9�O�>�۰�����o���-??���k�2W6;����4ǽc���DDB�S|!��`Ǩ����䘓���/n;/wQ��j��ܐϮ؇5t�"yZ���ҋ�}Í�·�A� ֔y�n�9'�k��#��j�Z�6������S{�x#QI�u�aBy�/�P�lN�pƻ�z3��M�L��g���4(SRT�oi�C�VpQ�)C8�D�b| 	:I^�v�HI�G���)�E��RDl&�[5I
��nŢ�Ă�#�:�nx�_������I��-�xiۘ�F*��J���E:�~����	�2�VȪ�]����a�+Yf s9{�g�����~�q��l�S�����~b=m�<�ߋ�Ώ$�D�x`��_*Ƌ��|��'�TuW�ݪo�m�{�81�EPS�b�
1FԎ�R {��ɇ�MB�
ٰzo��2�ǝ,Ί�X���\���@W�A����g#�R[�Q�w�F>	W���a�2�&�Iʳq+X�9d�@c���v��'
�M�#�Q6�)vm�°���<��I�Zx{�2!����S�����c!�8@�aee@�{i�].e�p��ƶ�hK�U�'�t-�0�Gq���@��@ۊ�E<י?x�18ŒY���$Q�f�����e��F�ϻW�#x�}��p]k�R�R?���7�Q����կ�������ka>$�Y#.�ҍ�|����v�(���I1Ͽ�/�P�S�=��5Mm��(�ŏv��or��b�ǽ����̴n� �;y[(� ���������磮+{���N�I�d��L��}��Zx�w�jK�^�k�+��F������8�WB�$B�p��[g��g7{��5��2Pg�=D-��At�E'%���l-&Z��S>.��e����#kЯ�7�f���@�e�+������6 �Ie���A���^+����D3�H�ӕ�� ��C%�\�i������o����a�m \�{`lR����	Z��"��N�L���)�-��Y�0�2,>Z�f2���x$��P���i#n��X�;��4~C��O9.�y�o��O+����,q3�ƾ��s����:��@�̳9ǄBV��ez'�?�t���r�&�B�#�eҢ��O@�7����p��G��TwUM�>}��g��2��%qOv���T�dS�+��됓!��B�y�	�"�
R�5d��`Bz'D��Y�W t]�v��� �
�8+։/37���G�v���Ю�`y�>����%}$��_i9������ˍ$<�S�,����ȫf�C��EO%9;}�l��Bb<��a�ߏ�FH,�������S�KC�����6o5w���czT<(5���)���Up�lO��ZB^P�i�����?�h	�z�b���*��.&��Z����9��Λ��yIu�0�r�ҡN�1�3�Q�)���f2�AK�}H�;�D����2:%0W:�+�~I8aߗP�lޝ����f�uɺ�`y�1�m�2lb�l
ȦP�`So�JQ>x��ωZ�Z8��X�/p�$�'t(e�W�os��oL��N�.�}9����Q�p��,N���J���DY��?7���⧁(��0��FEl�9y�W��	��N��M��U��ό�]d�q��q��ExiOX%^��_�z��ըM��z'�|C�{��_8uz�k�t����)���\ֳaVɩ�ۺb�E+s`90���o�A��6Tm���g���j��wI��	�*��~���Q �#Җ�a�=L� C��W�~!��#�FAh���|�K�����ȶ����j�7?ޛ�s�Ȥf�vb���<��6����Q�n$d�7�qQ�`jQ�U#]�	^�*Ӻvs����@���±U:�N�W���}m$�之�$�ɜ��y]�q$����3�ĝ�'QR
����U��O����WfW�F2�X�i�;n"��=��3z�HrW�~P���"l�+�jP����J#�{��'��F���K:����253�^	��p4i�[�<�Pt{��Q���C��t�hY�\|��h�u���aN?���zV�a�h:͡��>�&ȱ�P�X���}�=�g+�3#�`�5)ΌD����\9Q0�>�$n"���h���Vx\�B1ƽ�[�ͨ��Ri��/�by��+@�*f�@|����\�;��Q��~ۍ����R��݉�&c�y�,��$�G�e���<�S��#哞���� �Űf�ާy��x���o1��k2��=�|�=σ���]�@�o�r!��W]PRɧT\t+�ψx9+�O������X=��Z�5~�ξ�l~�Y�]h�NW`�:����Nb�ǒ&x¡�?�,�o׳)�����ߚ��n�	�Y��$�>m�Zys��YQ*'�W4L3R��wX8i��Δ�g#�S婰`H�Ѓv��r�H	�6m�Gȯ�`Px~UBʂ�������H!�XFe>y�⭨.� ��k(�(U��sv��gW�YG�-d��9"��$�������
*�.'^��*��]O�sE���g��'���;��,߇'��v.��'�`X�u85Z�}�칗'Yn��+��