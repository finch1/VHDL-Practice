--smi_int